`timescale 1ns/10ps
module huffman_DW01_add_0 ( A, B, CI, SUM, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [7:1] carry;

  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFXL U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  XOR3X1 U1_7 ( .A(A[7]), .B(B[7]), .C(carry[7]), .Y(SUM[7]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module huffman_DW01_add_1 ( A, B, CI, SUM, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [7:1] carry;

  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFXL U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  XOR3X1 U1_7 ( .A(A[7]), .B(B[7]), .C(carry[7]), .Y(SUM[7]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module huffman_DW01_add_2 ( A, B, CI, SUM, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [7:1] carry;

  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFXL U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  XOR3X1 U1_7 ( .A(A[7]), .B(B[7]), .C(carry[7]), .Y(SUM[7]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module huffman_DW01_add_3 ( A, B, CI, SUM, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [7:1] carry;

  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  XOR3X1 U1_7 ( .A(A[7]), .B(B[7]), .C(carry[7]), .Y(SUM[7]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module huffman_DW01_inc_0 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  ADDHXL U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  ADDHXL U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDHXL U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHXL U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHXL U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  ADDHXL U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  XOR2X1 U1 ( .A(carry[7]), .B(A[7]), .Y(SUM[7]) );
endmodule


module huffman_DW01_inc_1 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  ADDHXL U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  ADDHXL U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHXL U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHXL U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDHXL U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDHXL U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  CLKINVX1 U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1 U2 ( .A(carry[7]), .B(A[7]), .Y(SUM[7]) );
endmodule


module huffman_DW01_inc_2 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  ADDHXL U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  ADDHXL U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHXL U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDHXL U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHXL U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  ADDHXL U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  CLKINVX1 U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1 U2 ( .A(carry[7]), .B(A[7]), .Y(SUM[7]) );
endmodule


module huffman_DW01_inc_3 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  ADDHXL U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  ADDHXL U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHXL U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHXL U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDHXL U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDHXL U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  CLKINVX1 U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1 U2 ( .A(carry[7]), .B(A[7]), .Y(SUM[7]) );
endmodule


module huffman_DW01_inc_4 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  ADDHXL U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  ADDHXL U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDHXL U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHXL U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDHXL U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHXL U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  CLKINVX1 U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1 U2 ( .A(carry[7]), .B(A[7]), .Y(SUM[7]) );
endmodule


module huffman_DW01_inc_5 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  ADDHXL U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  ADDHXL U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHXL U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHXL U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDHXL U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDHXL U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  CLKINVX1 U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1 U2 ( .A(carry[7]), .B(A[7]), .Y(SUM[7]) );
endmodule


module huffman_DW01_inc_6 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  ADDHXL U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  ADDHXL U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDHXL U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHXL U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDHXL U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHXL U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  CLKINVX1 U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1 U2 ( .A(carry[7]), .B(A[7]), .Y(SUM[7]) );
endmodule


module huffman_DW01_inc_7 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  ADDHXL U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  ADDHXL U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHXL U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHXL U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDHXL U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDHXL U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  CLKINVX1 U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1 U2 ( .A(carry[7]), .B(A[7]), .Y(SUM[7]) );
endmodule


module huffman_DW01_inc_8 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  ADDHXL U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  ADDHXL U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDHXL U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHXL U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDHXL U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHXL U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  CLKINVX1 U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1 U2 ( .A(carry[7]), .B(A[7]), .Y(SUM[7]) );
endmodule


module huffman_DW01_inc_9 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  ADDHXL U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  ADDHXL U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHXL U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHXL U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDHXL U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDHXL U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  CLKINVX1 U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1 U2 ( .A(carry[7]), .B(A[7]), .Y(SUM[7]) );
endmodule


module huffman_DW01_inc_10 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  ADDHXL U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  ADDHXL U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  ADDHXL U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDHXL U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHXL U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHXL U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  XOR2X1 U1 ( .A(carry[7]), .B(A[7]), .Y(SUM[7]) );
endmodule


module huffman_DW01_inc_11 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  ADDHXL U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  ADDHXL U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHXL U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHXL U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDHXL U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDHXL U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  CLKINVX1 U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1 U2 ( .A(carry[7]), .B(A[7]), .Y(SUM[7]) );
endmodule


module huffman ( clk, reset, gray_valid, gray_data, CNT_valid, CNT1, CNT2, 
        CNT3, CNT4, CNT5, CNT6, code_valid, HC1, HC2, HC3, HC4, HC5, HC6, M1, 
        M2, M3, M4, M5, M6 );
  input [7:0] gray_data;
  output [7:0] CNT1;
  output [7:0] CNT2;
  output [7:0] CNT3;
  output [7:0] CNT4;
  output [7:0] CNT5;
  output [7:0] CNT6;
  output [7:0] HC1;
  output [7:0] HC2;
  output [7:0] HC3;
  output [7:0] HC4;
  output [7:0] HC5;
  output [7:0] HC6;
  output [7:0] M1;
  output [7:0] M2;
  output [7:0] M3;
  output [7:0] M4;
  output [7:0] M5;
  output [7:0] M6;
  input clk, reset, gray_valid;
  output CNT_valid, code_valid;
  wire   \symbol_value[0][7] , \symbol_value[0][6] , \symbol_value[0][5] ,
         \symbol_value[0][4] , \symbol_value[0][3] , \symbol_value[0][2] ,
         \symbol_value[0][1] , \symbol_value[0][0] , \symbol_value[1][7] ,
         \symbol_value[1][6] , \symbol_value[1][5] , \symbol_value[1][4] ,
         \symbol_value[1][3] , \symbol_value[1][2] , \symbol_value[1][1] ,
         \symbol_value[1][0] , \symbol_value[2][7] , \symbol_value[2][6] ,
         \symbol_value[2][5] , \symbol_value[2][4] , \symbol_value[2][3] ,
         \symbol_value[2][2] , \symbol_value[2][1] , \symbol_value[2][0] ,
         \symbol_value[3][7] , \symbol_value[3][6] , \symbol_value[3][5] ,
         \symbol_value[3][4] , \symbol_value[3][3] , \symbol_value[3][2] ,
         \symbol_value[3][1] , \symbol_value[3][0] , \symbol_value[4][7] ,
         \symbol_value[4][6] , \symbol_value[4][5] , \symbol_value[4][4] ,
         \symbol_value[4][3] , \symbol_value[4][2] , \symbol_value[4][1] ,
         \symbol_value[4][0] , \symbol_value[5][7] , \symbol_value[5][6] ,
         \symbol_value[5][5] , \symbol_value[5][4] , \symbol_value[5][3] ,
         \symbol_value[5][2] , \symbol_value[5][1] , \symbol_value[5][0] ,
         \symbol[3][5] , \symbol[3][4] , \symbol[3][3] , \symbol[3][2] ,
         \symbol[3][1] , \symbol[3][0] , \symbol[4][5] , \symbol[4][4] ,
         \symbol[4][3] , \symbol[4][2] , \symbol[4][1] , \symbol[4][0] ,
         \symbol[5][5] , \symbol[5][4] , \symbol[5][3] , \symbol[5][2] ,
         \symbol[5][1] , \symbol[5][0] , \C1[3][7] , \C1[3][6] , \C1[3][5] ,
         \C1[3][4] , \C1[3][3] , \C1[3][2] , \C1[3][1] , \C1[3][0] ,
         \C1[4][7] , \C1[4][6] , \C1[4][5] , \C1[4][4] , \C1[4][3] ,
         \C1[4][2] , \C1[4][1] , \C1[4][0] , \C2[2][7] , \C2[2][6] ,
         \C2[2][5] , \C2[2][4] , \C2[2][3] , \C2[2][2] , \C2[2][1] ,
         \C2[2][0] , \C2[3][7] , \C2[3][6] , \C2[3][5] , \C2[3][4] ,
         \C2[3][3] , \C2[3][2] , \C2[3][1] , \C2[3][0] , \C3[1][7] ,
         \C3[1][6] , \C3[1][5] , \C3[1][4] , \C3[1][3] , \C3[1][2] ,
         \C3[1][1] , \C3[1][0] , \C3[2][7] , \C3[2][6] , \C3[2][5] ,
         \C3[2][4] , \C3[2][3] , \C3[2][2] , \C3[2][1] , \C3[2][0] ,
         \C4[0][7] , \C4[0][5] , \C4[0][4] , \C4[0][3] , \C4[0][2] ,
         \C4[0][1] , \C4[0][0] , \C4[1][6] , \C4[1][4] , \C4[1][2] ,
         \C4[1][0] , N887, N888, N889, N890, N891, N892, N893, N894, N896,
         N897, N898, N899, N900, N901, N902, N903, N904, N905, N906, N907,
         N908, N909, N910, N911, N912, N913, N914, N915, N916, N917, N918,
         N919, N920, N921, N922, N923, N924, N925, N926, N927, N928, N929,
         N930, N931, N932, N933, N934, N935, N936, N937, N938, N939, N940,
         N941, N942, N943, N944, N945, N946, N947, N948, N949, N950, N951,
         N952, N953, N954, N955, N956, N957, N958, N959, N960, N961, N962,
         N963, N964, N965, N966, N967, N968, N969, N970, N971, N972, N973,
         N974, N976, N977, N978, N979, N980, N981, N982, N1143, N1144, N1145,
         N1146, N1147, N1148, N1149, N1150, N1726, N1727, N1728, N1729, N1730,
         N1731, N1732, N1733, N2254, N2255, N2256, N2257, N2258, N2259, N2260,
         N2261, N2775, N2776, N2777, N2778, N2779, N2780, N2781, N2782, N2784,
         n751, n752, n753, n754, n755, n756, n757, n758, n771, n772, n773,
         n774, n775, n776, n777, n778, n792, n793, n794, n795, n796, n797,
         n798, n799, n813, n814, n815, n816, n817, n818, n819, n820, n834,
         n835, n836, n837, n838, n839, n840, n841, n855, n856, n857, n858,
         n859, n860, n861, n862, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1019, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1042, n1043, n1044, n1045,
         n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
         n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
         n1066, n1067, n1068, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
         n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
         n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
         n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
         n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
         n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1126, n1127, n1128,
         n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
         n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
         n1149, n1150, n1151, n1152, n1154, n1155, n1156, n1157, n1158, n1159,
         n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
         n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
         n1180, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
         n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
         n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
         n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
         n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
         n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
         n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
         n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
         n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
         n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
         n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
         n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
         n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
         n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
         n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
         n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
         n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350,
         n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360,
         n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370,
         n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380,
         n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390,
         n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400,
         n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410,
         n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420,
         n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430,
         n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440,
         n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450,
         n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460,
         n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470,
         n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480,
         n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490,
         n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500,
         n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510,
         n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520,
         n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530,
         n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540,
         n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550,
         n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560,
         n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570,
         n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580,
         n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590,
         n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600,
         n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610,
         n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620,
         n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630,
         n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640,
         n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650,
         n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660,
         n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670,
         n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680,
         n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690,
         n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700,
         n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710,
         n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720,
         n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730,
         n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740,
         n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750,
         n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760,
         n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770,
         n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780,
         n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790,
         n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800,
         n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810,
         n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820,
         n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830,
         n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840,
         n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850,
         n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860,
         n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870,
         n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880,
         n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890,
         n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900,
         n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910,
         n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920,
         n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930,
         n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940,
         n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950,
         n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960,
         n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970,
         n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980,
         n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990,
         n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000,
         n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010,
         n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020,
         n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030,
         n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040,
         n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050,
         n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060,
         n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070,
         n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080,
         n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090,
         n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100,
         n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110,
         n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120,
         n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130,
         n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140,
         n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150,
         n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160,
         n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170,
         n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180,
         n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190,
         n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200,
         n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210,
         n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220,
         n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230,
         n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240,
         n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250,
         n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260,
         n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270,
         n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280,
         n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290,
         n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300,
         n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310,
         n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320,
         n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330,
         n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340,
         n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350,
         n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360,
         n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370,
         n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380,
         n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390,
         n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400,
         n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410,
         n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420,
         n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430,
         n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440,
         n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450,
         n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460,
         n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470,
         n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480,
         n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490,
         n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500,
         n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510,
         n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520,
         n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530,
         n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540,
         n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550,
         n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560,
         n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570,
         n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580,
         n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590,
         n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600,
         n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610,
         n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620,
         n2621, n2622, n2623, n2624, n2625;
  wire   [2:0] sort_stage;
  wire   [3:0] state;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1;

  huffman_DW01_add_0 add_587 ( .A({\C3[1][7] , \C3[1][6] , \C3[1][5] , 
        \C3[1][4] , \C3[1][3] , \C3[1][2] , \C3[1][1] , \C3[1][0] }), .B({
        \C3[2][7] , \C3[2][6] , \C3[2][5] , \C3[2][4] , \C3[2][3] , \C3[2][2] , 
        \C3[2][1] , \C3[2][0] }), .CI(1'b0), .SUM({N2782, N2781, N2780, N2779, 
        N2778, N2777, N2776, N2775}) );
  huffman_DW01_add_1 add_493 ( .A({\C2[2][7] , \C2[2][6] , \C2[2][5] , 
        \C2[2][4] , \C2[2][3] , \C2[2][2] , \C2[2][1] , \C2[2][0] }), .B({
        \C2[3][7] , \C2[3][6] , \C2[3][5] , \C2[3][4] , \C2[3][3] , \C2[3][2] , 
        \C2[3][1] , \C2[3][0] }), .CI(1'b0), .SUM({N2261, N2260, N2259, N2258, 
        N2257, N2256, N2255, N2254}) );
  huffman_DW01_add_2 add_386 ( .A({\C1[3][7] , \C1[3][6] , \C1[3][5] , 
        \C1[3][4] , \C1[3][3] , \C1[3][2] , \C1[3][1] , \C1[3][0] }), .B({
        \C1[4][7] , \C1[4][6] , \C1[4][5] , \C1[4][4] , \C1[4][3] , \C1[4][2] , 
        \C1[4][1] , \C1[4][0] }), .CI(1'b0), .SUM({N1733, N1732, N1731, N1730, 
        N1729, N1728, N1727, N1726}) );
  huffman_DW01_add_3 add_268 ( .A({\symbol_value[4][7] , \symbol_value[4][6] , 
        \symbol_value[4][5] , \symbol_value[4][4] , \symbol_value[4][3] , 
        \symbol_value[4][2] , \symbol_value[4][1] , \symbol_value[4][0] }), 
        .B({\symbol_value[5][7] , \symbol_value[5][6] , \symbol_value[5][5] , 
        \symbol_value[5][4] , \symbol_value[5][3] , \symbol_value[5][2] , 
        \symbol_value[5][1] , \symbol_value[5][0] }), .CI(1'b0), .SUM({N1150, 
        N1149, N1148, N1147, N1146, N1145, N1144, N1143}) );
  huffman_DW01_inc_0 add_133 ( .A({\symbol_value[5][7] , \symbol_value[5][6] , 
        \symbol_value[5][5] , \symbol_value[5][4] , \symbol_value[5][3] , 
        \symbol_value[5][2] , \symbol_value[5][1] , \symbol_value[5][0] }), 
        .SUM({N982, N981, N980, N979, N978, N977, N976, 
        SYNOPSYS_UNCONNECTED__0}) );
  huffman_DW01_inc_1 add_132 ( .A(CNT6), .SUM({N974, N973, N972, N971, N970, 
        N969, N968, N967}) );
  huffman_DW01_inc_2 add_129 ( .A({\symbol_value[4][7] , \symbol_value[4][6] , 
        \symbol_value[4][5] , \symbol_value[4][4] , \symbol_value[4][3] , 
        \symbol_value[4][2] , \symbol_value[4][1] , \symbol_value[4][0] }), 
        .SUM({N966, N965, N964, N963, N962, N961, N960, N959}) );
  huffman_DW01_inc_3 add_128 ( .A(CNT5), .SUM({N958, N957, N956, N955, N954, 
        N953, N952, N951}) );
  huffman_DW01_inc_4 add_125 ( .A({\symbol_value[3][7] , \symbol_value[3][6] , 
        \symbol_value[3][5] , \symbol_value[3][4] , \symbol_value[3][3] , 
        \symbol_value[3][2] , \symbol_value[3][1] , \symbol_value[3][0] }), 
        .SUM({N950, N949, N948, N947, N946, N945, N944, N943}) );
  huffman_DW01_inc_5 add_124 ( .A(CNT4), .SUM({N942, N941, N940, N939, N938, 
        N937, N936, N935}) );
  huffman_DW01_inc_6 add_121 ( .A({\symbol_value[2][7] , \symbol_value[2][6] , 
        \symbol_value[2][5] , \symbol_value[2][4] , \symbol_value[2][3] , 
        \symbol_value[2][2] , \symbol_value[2][1] , \symbol_value[2][0] }), 
        .SUM({N934, N933, N932, N931, N930, N929, N928, N927}) );
  huffman_DW01_inc_7 add_120 ( .A(CNT3), .SUM({N926, N925, N924, N923, N922, 
        N921, N920, N919}) );
  huffman_DW01_inc_8 add_117 ( .A({\symbol_value[1][7] , \symbol_value[1][6] , 
        \symbol_value[1][5] , \symbol_value[1][4] , \symbol_value[1][3] , 
        \symbol_value[1][2] , \symbol_value[1][1] , \symbol_value[1][0] }), 
        .SUM({N918, N917, N916, N915, N914, N913, N912, N911}) );
  huffman_DW01_inc_9 add_116 ( .A(CNT2), .SUM({N910, N909, N908, N907, N906, 
        N905, N904, N903}) );
  huffman_DW01_inc_10 add_113 ( .A({\symbol_value[0][7] , \symbol_value[0][6] , 
        \symbol_value[0][5] , \symbol_value[0][4] , \symbol_value[0][3] , 
        \symbol_value[0][2] , \symbol_value[0][1] , \symbol_value[0][0] }), 
        .SUM({N902, N901, N900, N899, N898, N897, N896, 
        SYNOPSYS_UNCONNECTED__1}) );
  huffman_DW01_inc_11 add_112 ( .A(CNT1), .SUM({N894, N893, N892, N891, N890, 
        N889, N888, N887}) );
  DFFRX1 CNT_valid_reg ( .D(n1418), .CK(clk), .RN(n2619), .Q(CNT_valid), .QN(
        n1017) );
  DFFRX1 \M6_reg[7]  ( .D(n1164), .CK(clk), .RN(n1743), .Q(M6[7]), .QN(n855)
         );
  DFFRX1 \M5_reg[7]  ( .D(n1136), .CK(clk), .RN(n1757), .Q(M5[7]), .QN(n834)
         );
  DFFRX1 \M4_reg[7]  ( .D(n1108), .CK(clk), .RN(n1754), .Q(M4[7]), .QN(n813)
         );
  DFFRX1 \M3_reg[7]  ( .D(n1080), .CK(clk), .RN(n1757), .Q(M3[7]), .QN(n792)
         );
  DFFRX1 \M2_reg[7]  ( .D(n1052), .CK(clk), .RN(n1752), .Q(M2[7]), .QN(n771)
         );
  DFFRX1 \M1_reg[7]  ( .D(n1032), .CK(clk), .RN(n1751), .Q(M1[7]), .QN(n751)
         );
  DFFRX1 \HC6_reg[3]  ( .D(n1179), .CK(clk), .RN(n1744), .Q(HC6[3]), .QN(n2509) );
  DFFRX1 \HC6_reg[2]  ( .D(n1178), .CK(clk), .RN(n1744), .Q(HC6[2]), .QN(n2510) );
  DFFRX1 \HC6_reg[1]  ( .D(n1177), .CK(clk), .RN(n1744), .Q(HC6[1]), .QN(n2512) );
  DFFRX1 \HC6_reg[0]  ( .D(n1176), .CK(clk), .RN(n1744), .Q(HC6[0]), .QN(n2514) );
  DFFRX1 \HC6_reg[7]  ( .D(n1175), .CK(clk), .RN(n1744), .Q(HC6[7]), .QN(n2505) );
  DFFRX1 \HC6_reg[6]  ( .D(n1174), .CK(clk), .RN(n1744), .Q(HC6[6]), .QN(n2506) );
  DFFRX1 \HC6_reg[5]  ( .D(n1173), .CK(clk), .RN(n1743), .Q(HC6[5]), .QN(n2507) );
  DFFRX1 \HC6_reg[4]  ( .D(n1172), .CK(clk), .RN(n1743), .Q(HC6[4]), .QN(n2508) );
  DFFRX1 \HC5_reg[3]  ( .D(n1151), .CK(clk), .RN(n1742), .Q(HC5[3]), .QN(n2519) );
  DFFRX1 \HC5_reg[2]  ( .D(n1150), .CK(clk), .RN(n1742), .Q(HC5[2]), .QN(n2520) );
  DFFRX1 \HC5_reg[1]  ( .D(n1149), .CK(clk), .RN(n1741), .Q(HC5[1]), .QN(n2522) );
  DFFRX1 \HC5_reg[7]  ( .D(n1147), .CK(clk), .RN(n1741), .Q(HC5[7]), .QN(n2516) );
  DFFRX1 \HC5_reg[6]  ( .D(n1146), .CK(clk), .RN(n1741), .Q(HC5[6]), .QN(n2517) );
  DFFRX1 \HC5_reg[5]  ( .D(n1145), .CK(clk), .RN(n1741), .Q(HC5[5]), .QN(n2518) );
  DFFRX1 \HC4_reg[3]  ( .D(n1123), .CK(clk), .RN(n1755), .Q(HC4[3]), .QN(n2528) );
  DFFRX1 \HC4_reg[2]  ( .D(n1122), .CK(clk), .RN(n1755), .Q(HC4[2]), .QN(n2529) );
  DFFRX1 \HC4_reg[1]  ( .D(n1121), .CK(clk), .RN(n1755), .Q(HC4[1]), .QN(n2531) );
  DFFRX1 \HC4_reg[7]  ( .D(n1119), .CK(clk), .RN(n1755), .Q(HC4[7]), .QN(n2525) );
  DFFRX1 \HC4_reg[6]  ( .D(n1118), .CK(clk), .RN(n1755), .Q(HC4[6]), .QN(n2526) );
  DFFRX1 \HC4_reg[5]  ( .D(n1117), .CK(clk), .RN(n1755), .Q(HC4[5]), .QN(n2527) );
  DFFRX1 \HC3_reg[3]  ( .D(n1095), .CK(clk), .RN(n1753), .Q(HC3[3]), .QN(n2537) );
  DFFRX1 \HC3_reg[2]  ( .D(n1094), .CK(clk), .RN(n1753), .Q(HC3[2]), .QN(n2538) );
  DFFRX1 \HC3_reg[1]  ( .D(n1093), .CK(clk), .RN(n1753), .Q(HC3[1]), .QN(n2540) );
  DFFRX1 \HC3_reg[7]  ( .D(n1091), .CK(clk), .RN(n1753), .Q(HC3[7]), .QN(n2534) );
  DFFRX1 \HC3_reg[6]  ( .D(n1090), .CK(clk), .RN(n1764), .Q(HC3[6]), .QN(n2535) );
  DFFRX1 \HC3_reg[5]  ( .D(n1089), .CK(clk), .RN(n1766), .Q(HC3[5]), .QN(n2536) );
  DFFRX1 \HC2_reg[3]  ( .D(n1067), .CK(clk), .RN(n1761), .Q(HC2[3]), .QN(n2546) );
  DFFRX1 \HC2_reg[2]  ( .D(n1066), .CK(clk), .RN(n1763), .Q(HC2[2]), .QN(n2547) );
  DFFRX1 \HC2_reg[1]  ( .D(n1065), .CK(clk), .RN(n1762), .Q(HC2[1]), .QN(n2549) );
  DFFRX1 \HC2_reg[7]  ( .D(n1063), .CK(clk), .RN(n1758), .Q(HC2[7]), .QN(n2543) );
  DFFRX1 \HC2_reg[6]  ( .D(n1062), .CK(clk), .RN(n1761), .Q(HC2[6]), .QN(n2544) );
  DFFRX1 \HC2_reg[5]  ( .D(n1061), .CK(clk), .RN(n1760), .Q(HC2[5]), .QN(n2545) );
  DFFRX1 \HC1_reg[7]  ( .D(n1031), .CK(clk), .RN(n1750), .Q(HC1[7]), .QN(n2552) );
  DFFRX1 \HC1_reg[6]  ( .D(n1030), .CK(clk), .RN(n1750), .Q(HC1[6]), .QN(n2553) );
  DFFRX1 \HC1_reg[5]  ( .D(n1029), .CK(clk), .RN(n1750), .Q(HC1[5]), .QN(n2554) );
  DFFRX1 \HC1_reg[3]  ( .D(n1027), .CK(clk), .RN(n1750), .Q(HC1[3]), .QN(n2555) );
  DFFRX1 \HC1_reg[2]  ( .D(n1026), .CK(clk), .RN(n1750), .Q(HC1[2]), .QN(n2556) );
  DFFRX1 \HC1_reg[1]  ( .D(n1025), .CK(clk), .RN(n1750), .Q(HC1[1]), .QN(n2558) );
  DFFRX1 code_valid_reg ( .D(n1424), .CK(clk), .RN(n1761), .Q(code_valid), 
        .QN(n1019) );
  DFFSX1 \symbol_reg[0][0]  ( .D(n1389), .CK(clk), .SN(n1756), .QN(n1651) );
  DFFSX1 \symbol_reg[1][1]  ( .D(n1384), .CK(clk), .SN(n1756), .QN(n1519) );
  DFFSX1 \symbol_reg[2][2]  ( .D(n1379), .CK(clk), .SN(n1756), .QN(n1485) );
  DFFRX1 \symbol_reg[2][0]  ( .D(n1391), .CK(clk), .RN(n1758), .QN(n1482) );
  DFFRX1 \symbol_reg[1][0]  ( .D(n1390), .CK(clk), .RN(n1750), .QN(n1520) );
  DFFRX1 \symbol_reg[2][1]  ( .D(n1385), .CK(clk), .RN(n1741), .QN(n1486) );
  DFFRX1 \symbol_reg[0][1]  ( .D(n1383), .CK(clk), .RN(n1757), .QN(n1650) );
  DFFRX1 \symbol_reg[1][2]  ( .D(n1378), .CK(clk), .RN(n1758), .QN(n1518) );
  DFFRX1 \symbol_reg[0][2]  ( .D(n1377), .CK(clk), .RN(n1748), .QN(n1649) );
  DFFRX1 \symbol_reg[2][3]  ( .D(n1373), .CK(clk), .RN(n1763), .QN(n1484) );
  DFFRX1 \symbol_reg[1][3]  ( .D(n1372), .CK(clk), .RN(n1751), .QN(n1517) );
  DFFRX1 \symbol_reg[0][3]  ( .D(n1371), .CK(clk), .RN(n1767), .QN(n1648) );
  DFFRX1 \symbol_reg[2][4]  ( .D(n1367), .CK(clk), .RN(n2619), .QN(n1483) );
  DFFRX1 \symbol_reg[1][4]  ( .D(n1366), .CK(clk), .RN(n1765), .QN(n1516) );
  DFFRX1 \symbol_reg[0][4]  ( .D(n1365), .CK(clk), .RN(n1762), .QN(n1647) );
  DFFRX1 \symbol_reg[2][5]  ( .D(n1361), .CK(clk), .RN(n1763), .QN(n1479) );
  DFFRX1 \symbol_reg[1][5]  ( .D(n1360), .CK(clk), .RN(n1756), .QN(n1487) );
  DFFRX1 \symbol_reg[0][5]  ( .D(n1359), .CK(clk), .RN(n1756), .QN(n1646) );
  DFFRX1 \C1_symbol_reg[1][5]  ( .D(n1291), .CK(clk), .RN(n1753), .QN(n1504)
         );
  DFFRX1 \C1_symbol_reg[0][5]  ( .D(n1290), .CK(clk), .RN(n1766), .QN(n1558)
         );
  DFFRX1 \C1_symbol_reg[1][4]  ( .D(n1286), .CK(clk), .RN(n1752), .QN(n1505)
         );
  DFFRX1 \C1_symbol_reg[0][4]  ( .D(n1285), .CK(clk), .RN(n1759), .QN(n1559)
         );
  DFFRX1 \C1_symbol_reg[1][3]  ( .D(n1281), .CK(clk), .RN(n1758), .QN(n1506)
         );
  DFFRX1 \C1_symbol_reg[0][3]  ( .D(n1280), .CK(clk), .RN(n1757), .QN(n1560)
         );
  DFFRX1 \C1_symbol_reg[1][2]  ( .D(n1276), .CK(clk), .RN(n1764), .QN(n1507)
         );
  DFFRX1 \C1_symbol_reg[0][2]  ( .D(n1275), .CK(clk), .RN(n1766), .QN(n1561)
         );
  DFFRX1 \C1_symbol_reg[1][1]  ( .D(n1271), .CK(clk), .RN(n1745), .QN(n1508)
         );
  DFFRX1 \C1_symbol_reg[0][1]  ( .D(n1270), .CK(clk), .RN(n1765), .QN(n1562)
         );
  DFFRX1 \C1_symbol_reg[1][0]  ( .D(n1266), .CK(clk), .RN(n1764), .QN(n1509)
         );
  DFFRX1 \C1_symbol_reg[0][0]  ( .D(n1265), .CK(clk), .RN(n1766), .QN(n1563)
         );
  DFFRX1 \C2_symbol_reg[1][5]  ( .D(n1189), .CK(clk), .RN(n1745), .QN(n1510)
         );
  DFFRX1 \C2_symbol_reg[0][5]  ( .D(n1188), .CK(clk), .RN(n1745), .QN(n1640)
         );
  DFFRX1 \C3_symbol_reg[0][5]  ( .D(n1185), .CK(clk), .RN(n1744), .QN(n1565)
         );
  DFFRX1 \C2_symbol_reg[1][4]  ( .D(n1161), .CK(clk), .RN(n1742), .QN(n1511)
         );
  DFFRX1 \C2_symbol_reg[0][4]  ( .D(n1160), .CK(clk), .RN(n1742), .QN(n1641)
         );
  DFFRX1 \C3_symbol_reg[0][4]  ( .D(n1157), .CK(clk), .RN(n1742), .QN(n1566)
         );
  DFFRX1 \C2_symbol_reg[1][3]  ( .D(n1133), .CK(clk), .RN(n1757), .QN(n1512)
         );
  DFFRX1 \C2_symbol_reg[0][3]  ( .D(n1132), .CK(clk), .RN(n1767), .QN(n1642)
         );
  DFFRX1 \C3_symbol_reg[0][3]  ( .D(n1129), .CK(clk), .RN(n1756), .QN(n1567)
         );
  DFFRX1 \C2_symbol_reg[1][2]  ( .D(n1105), .CK(clk), .RN(n1754), .QN(n1513)
         );
  DFFRX1 \C2_symbol_reg[0][2]  ( .D(n1104), .CK(clk), .RN(n1754), .QN(n1643)
         );
  DFFRX1 \C3_symbol_reg[0][2]  ( .D(n1101), .CK(clk), .RN(n1753), .QN(n1568)
         );
  DFFRX1 \C2_symbol_reg[1][1]  ( .D(n1077), .CK(clk), .RN(n1749), .QN(n1514)
         );
  DFFRX1 \C2_symbol_reg[0][1]  ( .D(n1076), .CK(clk), .RN(n1747), .QN(n1644)
         );
  DFFRX1 \C3_symbol_reg[0][1]  ( .D(n1073), .CK(clk), .RN(n1748), .QN(n1569)
         );
  DFFRX1 \C2_symbol_reg[1][0]  ( .D(n1049), .CK(clk), .RN(n1752), .QN(n1515)
         );
  DFFRX1 \C2_symbol_reg[0][0]  ( .D(n1048), .CK(clk), .RN(n1752), .QN(n1645)
         );
  DFFRX1 \C3_symbol_reg[0][0]  ( .D(n1045), .CK(clk), .RN(n1752), .QN(n1570)
         );
  DFFRX1 \HC5_reg[0]  ( .D(n1148), .CK(clk), .RN(n1741), .Q(HC5[0]) );
  DFFRX1 \HC5_reg[4]  ( .D(n1144), .CK(clk), .RN(n1741), .Q(HC5[4]) );
  DFFRX1 \HC4_reg[0]  ( .D(n1120), .CK(clk), .RN(n1755), .Q(HC4[0]) );
  DFFRX1 \HC4_reg[4]  ( .D(n1116), .CK(clk), .RN(n1755), .Q(HC4[4]) );
  DFFRX1 \HC3_reg[0]  ( .D(n1092), .CK(clk), .RN(n1753), .Q(HC3[0]) );
  DFFRX1 \HC3_reg[4]  ( .D(n1088), .CK(clk), .RN(n1767), .Q(HC3[4]) );
  DFFRX1 \HC2_reg[0]  ( .D(n1064), .CK(clk), .RN(n1765), .Q(HC2[0]) );
  DFFRX1 \HC2_reg[4]  ( .D(n1060), .CK(clk), .RN(n1757), .Q(HC2[4]) );
  DFFRX1 \HC1_reg[4]  ( .D(n1028), .CK(clk), .RN(n1750), .Q(HC1[4]) );
  DFFRX1 \HC1_reg[0]  ( .D(n1024), .CK(clk), .RN(n1755), .Q(HC1[0]) );
  DFFRX1 \M6_reg[1]  ( .D(n1170), .CK(clk), .RN(n1743), .Q(M6[1]), .QN(n861)
         );
  DFFRX1 \M6_reg[2]  ( .D(n1169), .CK(clk), .RN(n1743), .Q(M6[2]), .QN(n860)
         );
  DFFRX1 \M6_reg[3]  ( .D(n1168), .CK(clk), .RN(n1743), .Q(M6[3]), .QN(n859)
         );
  DFFRX1 \M6_reg[4]  ( .D(n1167), .CK(clk), .RN(n1743), .Q(M6[4]), .QN(n858)
         );
  DFFRX1 \M6_reg[5]  ( .D(n1166), .CK(clk), .RN(n1743), .Q(M6[5]), .QN(n857)
         );
  DFFRX1 \M6_reg[6]  ( .D(n1165), .CK(clk), .RN(n1743), .Q(M6[6]), .QN(n856)
         );
  DFFRX1 \M5_reg[1]  ( .D(n1142), .CK(clk), .RN(n1741), .Q(M5[1]), .QN(n840)
         );
  DFFRX1 \M5_reg[2]  ( .D(n1141), .CK(clk), .RN(n1741), .Q(M5[2]), .QN(n839)
         );
  DFFRX1 \M5_reg[3]  ( .D(n1140), .CK(clk), .RN(n1741), .Q(M5[3]), .QN(n838)
         );
  DFFRX1 \M5_reg[4]  ( .D(n1139), .CK(clk), .RN(n1741), .Q(M5[4]), .QN(n837)
         );
  DFFRX1 \M5_reg[5]  ( .D(n1138), .CK(clk), .RN(n1745), .Q(M5[5]), .QN(n836)
         );
  DFFRX1 \M5_reg[6]  ( .D(n1137), .CK(clk), .RN(n1763), .Q(M5[6]), .QN(n835)
         );
  DFFRX1 \M4_reg[1]  ( .D(n1114), .CK(clk), .RN(n1754), .Q(M4[1]), .QN(n819)
         );
  DFFRX1 \M4_reg[2]  ( .D(n1113), .CK(clk), .RN(n1754), .Q(M4[2]), .QN(n818)
         );
  DFFRX1 \M4_reg[3]  ( .D(n1112), .CK(clk), .RN(n1754), .Q(M4[3]), .QN(n817)
         );
  DFFRX1 \M4_reg[4]  ( .D(n1111), .CK(clk), .RN(n1754), .Q(M4[4]), .QN(n816)
         );
  DFFRX1 \M4_reg[5]  ( .D(n1110), .CK(clk), .RN(n1754), .Q(M4[5]), .QN(n815)
         );
  DFFRX1 \M4_reg[6]  ( .D(n1109), .CK(clk), .RN(n1754), .Q(M4[6]), .QN(n814)
         );
  DFFRX1 \M3_reg[1]  ( .D(n1086), .CK(clk), .RN(n1756), .Q(M3[1]), .QN(n798)
         );
  DFFRX1 \M3_reg[2]  ( .D(n1085), .CK(clk), .RN(n1749), .Q(M3[2]), .QN(n797)
         );
  DFFRX1 \M3_reg[3]  ( .D(n1084), .CK(clk), .RN(n1747), .Q(M3[3]), .QN(n796)
         );
  DFFRX1 \M3_reg[4]  ( .D(n1083), .CK(clk), .RN(n1755), .Q(M3[4]), .QN(n795)
         );
  DFFRX1 \M3_reg[5]  ( .D(n1082), .CK(clk), .RN(n1754), .Q(M3[5]), .QN(n794)
         );
  DFFRX1 \M3_reg[6]  ( .D(n1081), .CK(clk), .RN(n1747), .Q(M3[6]), .QN(n793)
         );
  DFFRX1 \M2_reg[1]  ( .D(n1058), .CK(clk), .RN(n1759), .Q(M2[1]), .QN(n777)
         );
  DFFRX1 \M2_reg[2]  ( .D(n1057), .CK(clk), .RN(n1764), .Q(M2[2]), .QN(n776)
         );
  DFFRX1 \M2_reg[3]  ( .D(n1056), .CK(clk), .RN(n1767), .Q(M2[3]), .QN(n775)
         );
  DFFRX1 \M2_reg[4]  ( .D(n1055), .CK(clk), .RN(n1752), .Q(M2[4]), .QN(n774)
         );
  DFFRX1 \M2_reg[5]  ( .D(n1054), .CK(clk), .RN(n1752), .Q(M2[5]), .QN(n773)
         );
  DFFRX1 \M2_reg[6]  ( .D(n1053), .CK(clk), .RN(n1752), .Q(M2[6]), .QN(n772)
         );
  DFFRX1 \M1_reg[1]  ( .D(n1038), .CK(clk), .RN(n1751), .Q(M1[1]), .QN(n757)
         );
  DFFRX1 \M1_reg[2]  ( .D(n1037), .CK(clk), .RN(n1751), .Q(M1[2]), .QN(n756)
         );
  DFFRX1 \M1_reg[3]  ( .D(n1036), .CK(clk), .RN(n1751), .Q(M1[3]), .QN(n755)
         );
  DFFRX1 \M1_reg[4]  ( .D(n1035), .CK(clk), .RN(n1751), .Q(M1[4]), .QN(n754)
         );
  DFFRX1 \M1_reg[5]  ( .D(n1034), .CK(clk), .RN(n1751), .Q(M1[5]), .QN(n753)
         );
  DFFRX1 \M1_reg[6]  ( .D(n1033), .CK(clk), .RN(n1751), .Q(M1[6]), .QN(n752)
         );
  DFFRX1 \symbol_reg[3][0]  ( .D(n1394), .CK(clk), .RN(n1764), .Q(
        \symbol[3][0] ), .QN(n1553) );
  DFFRX1 \symbol_reg[3][1]  ( .D(n1388), .CK(clk), .RN(n1749), .Q(
        \symbol[3][1] ), .QN(n1554) );
  DFFRX1 \symbol_reg[3][2]  ( .D(n1382), .CK(clk), .RN(n1763), .Q(
        \symbol[3][2] ), .QN(n1555) );
  DFFRX1 \symbol_reg[3][4]  ( .D(n1370), .CK(clk), .RN(n1742), .Q(
        \symbol[3][4] ), .QN(n1556) );
  DFFRX1 \symbol_reg[3][5]  ( .D(n1364), .CK(clk), .RN(n1749), .Q(
        \symbol[3][5] ), .QN(n1522) );
  DFFRX1 \M6_reg[0]  ( .D(n1171), .CK(clk), .RN(n1743), .Q(M6[0]), .QN(n862)
         );
  DFFRX1 \M5_reg[0]  ( .D(n1143), .CK(clk), .RN(n1741), .Q(M5[0]), .QN(n841)
         );
  DFFRX1 \M4_reg[0]  ( .D(n1115), .CK(clk), .RN(n1755), .Q(M4[0]), .QN(n820)
         );
  DFFRX1 \M3_reg[0]  ( .D(n1087), .CK(clk), .RN(n1743), .Q(M3[0]), .QN(n799)
         );
  DFFRX1 \M2_reg[0]  ( .D(n1059), .CK(clk), .RN(n1766), .Q(M2[0]), .QN(n778)
         );
  DFFRX1 \M1_reg[0]  ( .D(n1039), .CK(clk), .RN(n1751), .Q(M1[0]), .QN(n758)
         );
  DFFSX1 \symbol_reg[3][3]  ( .D(n1376), .CK(clk), .SN(n1756), .Q(
        \symbol[3][3] ), .QN(n1557) );
  DFFRX1 \CNT6_reg[7]  ( .D(n1470), .CK(clk), .RN(n1757), .Q(CNT6[7]) );
  DFFRX1 \CNT4_reg[7]  ( .D(n1462), .CK(clk), .RN(n1762), .Q(CNT4[7]) );
  DFFRX1 \CNT2_reg[7]  ( .D(n1454), .CK(clk), .RN(n1758), .Q(CNT2[7]) );
  DFFRX1 \CNT5_reg[7]  ( .D(n1446), .CK(clk), .RN(n1753), .Q(CNT5[7]) );
  DFFRX1 \CNT3_reg[7]  ( .D(n1438), .CK(clk), .RN(n1767), .Q(CNT3[7]) );
  DFFRX1 \CNT1_reg[7]  ( .D(n1430), .CK(clk), .RN(n1759), .Q(CNT1[7]) );
  DFFRX1 \C1_symbol_reg[2][5]  ( .D(n1292), .CK(clk), .RN(n1765), .Q(n2612) );
  DFFRX1 \C1_symbol_reg[2][4]  ( .D(n1287), .CK(clk), .RN(n1763), .Q(n2613) );
  DFFRX1 \C1_symbol_reg[2][3]  ( .D(n1282), .CK(clk), .RN(n1767), .Q(n2614) );
  DFFRX1 \C1_symbol_reg[2][2]  ( .D(n1277), .CK(clk), .RN(n1756), .Q(n2615) );
  DFFRX1 \C1_symbol_reg[2][1]  ( .D(n1272), .CK(clk), .RN(n1758), .Q(n2616) );
  DFFRX1 \C1_symbol_reg[2][0]  ( .D(n1267), .CK(clk), .RN(n1758), .Q(n2617) );
  DFFRX1 \CNT6_reg[2]  ( .D(n1475), .CK(clk), .RN(n1752), .Q(CNT6[2]) );
  DFFRX1 \CNT6_reg[3]  ( .D(n1474), .CK(clk), .RN(n1759), .Q(CNT6[3]) );
  DFFRX1 \CNT6_reg[4]  ( .D(n1473), .CK(clk), .RN(n1758), .Q(CNT6[4]) );
  DFFRX1 \CNT6_reg[5]  ( .D(n1472), .CK(clk), .RN(n1761), .Q(CNT6[5]) );
  DFFRX1 \CNT6_reg[6]  ( .D(n1471), .CK(clk), .RN(n1760), .Q(CNT6[6]) );
  DFFRX1 \CNT4_reg[2]  ( .D(n1467), .CK(clk), .RN(n2619), .Q(CNT4[2]) );
  DFFRX1 \CNT4_reg[3]  ( .D(n1466), .CK(clk), .RN(n1761), .Q(CNT4[3]) );
  DFFRX1 \CNT4_reg[4]  ( .D(n1465), .CK(clk), .RN(n1764), .Q(CNT4[4]) );
  DFFRX1 \CNT4_reg[5]  ( .D(n1464), .CK(clk), .RN(n1760), .Q(CNT4[5]) );
  DFFRX1 \CNT4_reg[6]  ( .D(n1463), .CK(clk), .RN(n1763), .Q(CNT4[6]) );
  DFFRX1 \CNT2_reg[2]  ( .D(n1459), .CK(clk), .RN(n1762), .Q(CNT2[2]) );
  DFFRX1 \CNT2_reg[3]  ( .D(n1458), .CK(clk), .RN(n1754), .Q(CNT2[3]) );
  DFFRX1 \CNT2_reg[4]  ( .D(n1457), .CK(clk), .RN(n1743), .Q(CNT2[4]) );
  DFFRX1 \CNT2_reg[5]  ( .D(n1456), .CK(clk), .RN(n1765), .Q(CNT2[5]) );
  DFFRX1 \CNT2_reg[6]  ( .D(n1455), .CK(clk), .RN(n1764), .Q(CNT2[6]) );
  DFFRX1 \CNT5_reg[2]  ( .D(n1451), .CK(clk), .RN(n1766), .Q(CNT5[2]) );
  DFFRX1 \CNT5_reg[3]  ( .D(n1450), .CK(clk), .RN(n1765), .Q(CNT5[3]) );
  DFFRX1 \CNT5_reg[4]  ( .D(n1449), .CK(clk), .RN(n1764), .Q(CNT5[4]) );
  DFFRX1 \CNT5_reg[5]  ( .D(n1448), .CK(clk), .RN(n1766), .Q(CNT5[5]) );
  DFFRX1 \CNT5_reg[6]  ( .D(n1447), .CK(clk), .RN(n1757), .Q(CNT5[6]) );
  DFFRX1 \CNT3_reg[2]  ( .D(n1443), .CK(clk), .RN(n1753), .Q(CNT3[2]) );
  DFFRX1 \CNT3_reg[3]  ( .D(n1442), .CK(clk), .RN(n1758), .Q(CNT3[3]) );
  DFFRX1 \CNT3_reg[4]  ( .D(n1441), .CK(clk), .RN(n1765), .Q(CNT3[4]) );
  DFFRX1 \CNT3_reg[5]  ( .D(n1440), .CK(clk), .RN(n1767), .Q(CNT3[5]) );
  DFFRX1 \CNT3_reg[6]  ( .D(n1439), .CK(clk), .RN(n1759), .Q(CNT3[6]) );
  DFFRX1 \CNT1_reg[2]  ( .D(n1435), .CK(clk), .RN(n1765), .Q(CNT1[2]) );
  DFFRX1 \CNT1_reg[3]  ( .D(n1434), .CK(clk), .RN(n1763), .Q(CNT1[3]) );
  DFFRX1 \CNT1_reg[4]  ( .D(n1433), .CK(clk), .RN(n1761), .Q(CNT1[4]) );
  DFFRX1 \CNT1_reg[5]  ( .D(n1432), .CK(clk), .RN(n1760), .Q(CNT1[5]) );
  DFFRX1 \CNT1_reg[6]  ( .D(n1431), .CK(clk), .RN(n1763), .Q(CNT1[6]) );
  DFFRX1 \HC_length_reg[5][2]  ( .D(n1180), .CK(clk), .RN(n1744), .Q(n2515), 
        .QN(n1637) );
  DFFRX1 \HC_length_reg[5][1]  ( .D(n2625), .CK(clk), .RN(n1744), .Q(n2511), 
        .QN(n1638) );
  DFFRX1 \HC_length_reg[5][0]  ( .D(n1182), .CK(clk), .RN(n1744), .Q(n2513), 
        .QN(n1552) );
  DFFRX1 \CNT6_reg[1]  ( .D(n1476), .CK(clk), .RN(n1753), .Q(CNT6[1]) );
  DFFRX1 \CNT4_reg[1]  ( .D(n1468), .CK(clk), .RN(n1762), .Q(CNT4[1]) );
  DFFRX1 \CNT2_reg[1]  ( .D(n1460), .CK(clk), .RN(n1759), .Q(CNT2[1]) );
  DFFRX1 \CNT5_reg[1]  ( .D(n1452), .CK(clk), .RN(n1767), .Q(CNT5[1]) );
  DFFRX1 \CNT3_reg[1]  ( .D(n1444), .CK(clk), .RN(n1763), .Q(CNT3[1]) );
  DFFRX1 \CNT1_reg[1]  ( .D(n1436), .CK(clk), .RN(n1762), .Q(CNT1[1]) );
  DFFRX1 \C1_reg[0][7]  ( .D(n1328), .CK(clk), .RN(n1757), .QN(n1009) );
  DFFRX1 \C2_reg[0][7]  ( .D(n1259), .CK(clk), .RN(n1741), .QN(n940) );
  DFFRX1 \CNT6_reg[0]  ( .D(n1477), .CK(clk), .RN(n1741), .Q(CNT6[0]) );
  DFFRX1 \CNT4_reg[0]  ( .D(n1469), .CK(clk), .RN(n1761), .Q(CNT4[0]) );
  DFFRX1 \CNT2_reg[0]  ( .D(n1461), .CK(clk), .RN(n1767), .Q(CNT2[0]) );
  DFFRX1 \CNT5_reg[0]  ( .D(n1453), .CK(clk), .RN(n1766), .Q(CNT5[0]) );
  DFFRX1 \CNT3_reg[0]  ( .D(n1445), .CK(clk), .RN(n1757), .Q(CNT3[0]) );
  DFFRX1 \CNT1_reg[0]  ( .D(n1437), .CK(clk), .RN(n1761), .Q(CNT1[0]) );
  DFFRX1 \HC_length_reg[4][0]  ( .D(n1154), .CK(clk), .RN(n1742), .Q(n2523), 
        .QN(n1627) );
  DFFRX1 \HC_length_reg[3][0]  ( .D(n1126), .CK(clk), .RN(n1755), .Q(n2532), 
        .QN(n1628) );
  DFFRX1 \HC_length_reg[2][0]  ( .D(n1098), .CK(clk), .RN(n1753), .Q(n2541), 
        .QN(n1629) );
  DFFRX1 \HC_length_reg[1][0]  ( .D(n1070), .CK(clk), .RN(n1752), .Q(n2550), 
        .QN(n1630) );
  DFFRX1 \HC_length_reg[0][0]  ( .D(n1042), .CK(clk), .RN(n1751), .Q(n2559), 
        .QN(n1631) );
  DFFRX1 \HC_length_reg[4][1]  ( .D(n2624), .CK(clk), .RN(n1742), .Q(n2521) );
  DFFRX1 \HC_length_reg[3][1]  ( .D(n2623), .CK(clk), .RN(n1755), .Q(n2530) );
  DFFRX1 \HC_length_reg[2][1]  ( .D(n2622), .CK(clk), .RN(n1753), .Q(n2539) );
  DFFRX1 \HC_length_reg[1][1]  ( .D(n2621), .CK(clk), .RN(n1751), .Q(n2548) );
  DFFRX1 \HC_length_reg[0][1]  ( .D(n2620), .CK(clk), .RN(n1751), .Q(n2557) );
  DFFRX1 \C4_reg[1][7]  ( .D(n1206), .CK(clk), .RN(n1746), .QN(n889) );
  DFFRX1 \C4_reg[0][7]  ( .D(n1207), .CK(clk), .RN(n1746), .Q(\C4[0][7] ), 
        .QN(n890) );
  DFFSX1 \symbol_reg[5][5]  ( .D(n1362), .CK(clk), .SN(n1756), .Q(
        \symbol[5][5] ), .QN(n1684) );
  DFFRX1 \C4_reg[1][6]  ( .D(n1192), .CK(clk), .RN(n1745), .Q(\C4[1][6] ), 
        .QN(n875) );
  DFFRX1 \HC_length_reg[4][2]  ( .D(n1152), .CK(clk), .RN(n1742), .Q(n2524), 
        .QN(n1632) );
  DFFRX1 \HC_length_reg[3][2]  ( .D(n1124), .CK(clk), .RN(n1755), .Q(n2533), 
        .QN(n1633) );
  DFFRX1 \HC_length_reg[2][2]  ( .D(n1096), .CK(clk), .RN(n1753), .Q(n2542), 
        .QN(n1634) );
  DFFRX1 \HC_length_reg[1][2]  ( .D(n1068), .CK(clk), .RN(n1741), .Q(n2551), 
        .QN(n1635) );
  DFFRX1 \HC_length_reg[0][2]  ( .D(n1040), .CK(clk), .RN(n1751), .Q(n2560), 
        .QN(n1636) );
  DFFRX1 \C1_reg[4][4]  ( .D(n1310), .CK(clk), .RN(n1757), .Q(\C1[4][4] ), 
        .QN(n992) );
  DFFRX1 \C1_reg[4][2]  ( .D(n1300), .CK(clk), .RN(n1765), .Q(\C1[4][2] ), 
        .QN(n982) );
  DFFRX1 \C1_reg[4][0]  ( .D(n1332), .CK(clk), .RN(n1750), .Q(\C1[4][0] ), 
        .QN(n1015) );
  DFFRX1 \C2_reg[3][7]  ( .D(n1232), .CK(clk), .RN(n1748), .Q(\C2[3][7] ), 
        .QN(n942) );
  DFFRX1 \C1_reg[4][7]  ( .D(n1294), .CK(clk), .RN(n1762), .Q(\C1[4][7] ), 
        .QN(n1012) );
  DFFRX1 \C3_reg[2][7]  ( .D(n1231), .CK(clk), .RN(n1748), .Q(\C3[2][7] ), 
        .QN(n914) );
  DFFRX1 \C1_reg[0][0]  ( .D(n1326), .CK(clk), .RN(n1761), .Q(n1602), .QN(
        n1007) );
  DFFRX1 \C2_reg[0][6]  ( .D(n1255), .CK(clk), .RN(n1742), .Q(n1595), .QN(n935) );
  DFFRX1 \C2_reg[0][0]  ( .D(n1233), .CK(clk), .RN(n1749), .Q(n1603), .QN(n939) );
  DFFRX1 \C3_reg[2][6]  ( .D(n1210), .CK(clk), .RN(n1747), .Q(\C3[2][6] ), 
        .QN(n893) );
  DFFRX1 \C1_reg[4][1]  ( .D(n1295), .CK(clk), .RN(n1760), .Q(\C1[4][1] ), 
        .QN(n977) );
  DFFRX1 \C3_reg[0][6]  ( .D(n1208), .CK(clk), .RN(n1746), .Q(n1599), .QN(n891) );
  DFFRX1 \C1_reg[0][6]  ( .D(n1322), .CK(clk), .RN(n1763), .Q(n1598), .QN(
        n1003) );
  DFFRX1 \C3_reg[0][3]  ( .D(n1217), .CK(clk), .RN(n1747), .QN(n900) );
  DFFRX1 \C2_reg[2][7]  ( .D(n1261), .CK(clk), .RN(n1746), .Q(\C2[2][7] ), 
        .QN(n943) );
  DFFRX1 \C1_reg[0][3]  ( .D(n1307), .CK(clk), .RN(n1763), .QN(n988) );
  DFFRX1 \C2_reg[0][3]  ( .D(n1243), .CK(clk), .RN(n1749), .QN(n923) );
  DFFRX1 \C1_reg[4][3]  ( .D(n1305), .CK(clk), .RN(n1762), .Q(\C1[4][3] ), 
        .QN(n987) );
  DFFRX1 \C2_reg[0][4]  ( .D(n1247), .CK(clk), .RN(n1750), .QN(n927) );
  DFFRX1 \C3_reg[0][2]  ( .D(n1220), .CK(clk), .RN(n1747), .QN(n903) );
  DFFRX1 \C3_reg[1][7]  ( .D(n1230), .CK(clk), .RN(n1748), .Q(\C3[1][7] ), 
        .QN(n913) );
  DFFRX1 \C1_reg[0][4]  ( .D(n1312), .CK(clk), .RN(n1756), .QN(n993) );
  DFFRX1 \C1_reg[4][6]  ( .D(n1320), .CK(clk), .RN(n1764), .Q(\C1[4][6] ), 
        .QN(n1002) );
  DFFRX1 \C1_reg[0][2]  ( .D(n1302), .CK(clk), .RN(n1760), .QN(n983) );
  DFFRX1 \C2_reg[0][2]  ( .D(n1239), .CK(clk), .RN(n1749), .QN(n919) );
  DFFRX1 \C3_reg[0][7]  ( .D(n1229), .CK(clk), .RN(n1748), .QN(n912) );
  DFFRX1 \C2_reg[1][7]  ( .D(n1260), .CK(clk), .RN(n1745), .Q(n1607), .QN(n941) );
  DFFRX1 \C4_reg[0][0]  ( .D(n1205), .CK(clk), .RN(n1746), .Q(\C4[0][0] ), 
        .QN(n888) );
  DFFRX1 \C4_reg[1][0]  ( .D(n1204), .CK(clk), .RN(n1746), .Q(\C4[1][0] ), 
        .QN(n887) );
  DFFRX1 \C4_reg[1][1]  ( .D(n1202), .CK(clk), .RN(n1746), .QN(n885) );
  DFFRX1 \C4_reg[1][3]  ( .D(n1198), .CK(clk), .RN(n1746), .QN(n881) );
  DFFRX1 \C4_reg[1][5]  ( .D(n1194), .CK(clk), .RN(n1745), .QN(n877) );
  DFFRX1 \C4_reg[0][6]  ( .D(n1193), .CK(clk), .RN(n1745), .QN(n876) );
  DFFRX1 \C4_symbol_reg[0][5]  ( .D(n1183), .CK(clk), .RN(n1744), .Q(n2561), 
        .QN(n1678) );
  DFFRX1 \C4_symbol_reg[0][4]  ( .D(n1155), .CK(clk), .RN(n1742), .Q(n2563), 
        .QN(n1679) );
  DFFRX1 \C4_symbol_reg[0][3]  ( .D(n1127), .CK(clk), .RN(n1757), .Q(n2565), 
        .QN(n1680) );
  DFFRX1 \C4_symbol_reg[0][2]  ( .D(n1099), .CK(clk), .RN(n1753), .Q(n2567), 
        .QN(n1681) );
  DFFRX1 \C4_symbol_reg[0][1]  ( .D(n1071), .CK(clk), .RN(n1742), .Q(n2569), 
        .QN(n1682) );
  DFFRX1 \C4_symbol_reg[0][0]  ( .D(n1043), .CK(clk), .RN(n1751), .Q(n2571), 
        .QN(n1683) );
  DFFRX1 \C4_symbol_reg[1][5]  ( .D(n1184), .CK(clk), .RN(n1744), .Q(n2562), 
        .QN(n1503) );
  DFFRX1 \C4_symbol_reg[1][4]  ( .D(n1156), .CK(clk), .RN(n1742), .Q(n2564), 
        .QN(n1488) );
  DFFRX1 \C4_symbol_reg[1][3]  ( .D(n1128), .CK(clk), .RN(n1766), .Q(n2566), 
        .QN(n1489) );
  DFFRX1 \C4_symbol_reg[1][2]  ( .D(n1100), .CK(clk), .RN(n1753), .Q(n2568), 
        .QN(n1490) );
  DFFRX1 \C4_symbol_reg[1][1]  ( .D(n1072), .CK(clk), .RN(n1746), .Q(n2570), 
        .QN(n1491) );
  DFFRX1 \C4_symbol_reg[1][0]  ( .D(n1044), .CK(clk), .RN(n1752), .Q(n2572), 
        .QN(n1492) );
  DFFRX1 \C4_reg[0][1]  ( .D(n1203), .CK(clk), .RN(n1746), .Q(\C4[0][1] ), 
        .QN(n886) );
  DFFRX1 \symbol_reg[4][5]  ( .D(n1363), .CK(clk), .RN(n1763), .Q(
        \symbol[4][5] ), .QN(n1564) );
  DFFRX1 \C1_symbol_reg[4][5]  ( .D(n1289), .CK(clk), .RN(n1759), .Q(n2600), 
        .QN(n1671) );
  DFFRX1 \C1_symbol_reg[4][4]  ( .D(n1284), .CK(clk), .RN(n1756), .Q(n2601), 
        .QN(n1666) );
  DFFRX1 \C1_symbol_reg[4][3]  ( .D(n1279), .CK(clk), .RN(n1748), .Q(n2602), 
        .QN(n1667) );
  DFFRX1 \C1_symbol_reg[4][2]  ( .D(n1274), .CK(clk), .RN(n1761), .Q(n2603), 
        .QN(n1668) );
  DFFRX1 \C1_symbol_reg[4][1]  ( .D(n1269), .CK(clk), .RN(n1744), .Q(n2604), 
        .QN(n1669) );
  DFFRX1 \C1_symbol_reg[4][0]  ( .D(n1264), .CK(clk), .RN(n1750), .Q(n2605), 
        .QN(n1670) );
  DFFRX1 \C2_symbol_reg[3][5]  ( .D(n1191), .CK(clk), .RN(n1745), .Q(n2587), 
        .QN(n1546) );
  DFFRX1 \C3_symbol_reg[2][5]  ( .D(n1187), .CK(clk), .RN(n1745), .Q(n2574), 
        .QN(n1672) );
  DFFRX1 \C2_symbol_reg[3][4]  ( .D(n1163), .CK(clk), .RN(n1743), .Q(n2588), 
        .QN(n1547) );
  DFFRX1 \C3_symbol_reg[2][4]  ( .D(n1159), .CK(clk), .RN(n1742), .Q(n2575), 
        .QN(n1673) );
  DFFRX1 \C2_symbol_reg[3][3]  ( .D(n1135), .CK(clk), .RN(n1764), .Q(n2589), 
        .QN(n1548) );
  DFFRX1 \C3_symbol_reg[2][3]  ( .D(n1131), .CK(clk), .RN(n1766), .Q(n2576), 
        .QN(n1674) );
  DFFRX1 \C2_symbol_reg[3][2]  ( .D(n1107), .CK(clk), .RN(n1754), .Q(n2590), 
        .QN(n1549) );
  DFFRX1 \C3_symbol_reg[2][2]  ( .D(n1103), .CK(clk), .RN(n1754), .Q(n2577), 
        .QN(n1675) );
  DFFRX1 \C2_symbol_reg[3][1]  ( .D(n1079), .CK(clk), .RN(n1745), .Q(n2591), 
        .QN(n1550) );
  DFFRX1 \C3_symbol_reg[2][1]  ( .D(n1075), .CK(clk), .RN(n1743), .Q(n2578), 
        .QN(n1676) );
  DFFRX1 \C2_symbol_reg[3][0]  ( .D(n1051), .CK(clk), .RN(n1752), .Q(n2592), 
        .QN(n1551) );
  DFFRX1 \C3_symbol_reg[2][0]  ( .D(n1047), .CK(clk), .RN(n1752), .Q(n2579), 
        .QN(n1677) );
  DFFRX1 \C4_reg[0][3]  ( .D(n1199), .CK(clk), .RN(n1746), .Q(\C4[0][3] ), 
        .QN(n882) );
  DFFRX1 \C2_reg[3][4]  ( .D(n1246), .CK(clk), .RN(n1750), .Q(\C2[3][4] ), 
        .QN(n929) );
  DFFRX1 \C3_symbol_reg[1][5]  ( .D(n1186), .CK(clk), .RN(n1745), .Q(n2580), 
        .QN(n1497) );
  DFFRX1 \C3_symbol_reg[1][4]  ( .D(n1158), .CK(clk), .RN(n1742), .Q(n2581), 
        .QN(n1498) );
  DFFRX1 \C3_symbol_reg[1][3]  ( .D(n1130), .CK(clk), .RN(n1759), .Q(n2582), 
        .QN(n1499) );
  DFFRX1 \C3_symbol_reg[1][2]  ( .D(n1102), .CK(clk), .RN(n1753), .Q(n2583), 
        .QN(n1500) );
  DFFRX1 \C3_symbol_reg[1][1]  ( .D(n1074), .CK(clk), .RN(n1744), .Q(n2584), 
        .QN(n1501) );
  DFFRX1 \C3_symbol_reg[1][0]  ( .D(n1046), .CK(clk), .RN(n1752), .Q(n2585), 
        .QN(n1502) );
  DFFRX1 \C2_reg[3][0]  ( .D(n1262), .CK(clk), .RN(n1760), .Q(\C2[3][0] ), 
        .QN(n945) );
  DFFRX1 \C3_reg[2][2]  ( .D(n1222), .CK(clk), .RN(n1748), .Q(\C3[2][2] ), 
        .QN(n905) );
  DFFRX1 \C2_symbol_reg[2][5]  ( .D(n1190), .CK(clk), .RN(n1745), .Q(n2593), 
        .QN(n1660) );
  DFFRX1 \C2_symbol_reg[2][4]  ( .D(n1162), .CK(clk), .RN(n1743), .Q(n2594), 
        .QN(n1661) );
  DFFRX1 \C2_symbol_reg[2][3]  ( .D(n1134), .CK(clk), .RN(n1746), .Q(n2595), 
        .QN(n1662) );
  DFFRX1 \C2_symbol_reg[2][2]  ( .D(n1106), .CK(clk), .RN(n1754), .Q(n2596), 
        .QN(n1663) );
  DFFRX1 \C2_symbol_reg[2][1]  ( .D(n1078), .CK(clk), .RN(n1755), .Q(n2597), 
        .QN(n1664) );
  DFFRX1 \C2_symbol_reg[2][0]  ( .D(n1050), .CK(clk), .RN(n1752), .Q(n2598), 
        .QN(n1665) );
  DFFRX1 \C3_reg[2][0]  ( .D(n1226), .CK(clk), .RN(n1748), .Q(\C3[2][0] ), 
        .QN(n910) );
  DFFRX1 \C2_reg[2][6]  ( .D(n1257), .CK(clk), .RN(n1743), .Q(\C2[2][6] ), 
        .QN(n938) );
  DFFRX1 \C3_reg[1][0]  ( .D(n1228), .CK(clk), .RN(n1748), .Q(\C3[1][0] ), 
        .QN(n911) );
  DFFRX1 \C3_reg[1][1]  ( .D(n1224), .CK(clk), .RN(n1748), .Q(\C3[1][1] ), 
        .QN(n907) );
  DFFRX1 \C3_reg[1][4]  ( .D(n1215), .CK(clk), .RN(n1747), .Q(\C3[1][4] ), 
        .QN(n898) );
  DFFRX1 \C2_reg[3][5]  ( .D(n1250), .CK(clk), .RN(n1750), .Q(\C2[3][5] ), 
        .QN(n933) );
  DFFRX1 \C1_reg[0][1]  ( .D(n1297), .CK(clk), .RN(n1764), .Q(n1536), .QN(n978) );
  DFFRX1 \C2_reg[0][1]  ( .D(n1235), .CK(clk), .RN(n1749), .Q(n1537), .QN(n915) );
  DFFRX1 \C3_reg[0][0]  ( .D(n1227), .CK(clk), .RN(n1748), .QN(n909) );
  DFFRX1 \C1_reg[4][5]  ( .D(n1315), .CK(clk), .RN(n1752), .Q(\C1[4][5] ), 
        .QN(n997) );
  DFFRX1 \C2_reg[3][1]  ( .D(n1234), .CK(clk), .RN(n1749), .Q(\C2[3][1] ), 
        .QN(n917) );
  DFFRX1 \C1_symbol_reg[3][5]  ( .D(n1293), .CK(clk), .RN(n1766), .Q(n2606), 
        .QN(n1576) );
  DFFRX1 \C1_symbol_reg[3][4]  ( .D(n1288), .CK(clk), .RN(n1767), .Q(n2607), 
        .QN(n1573) );
  DFFRX1 \C1_symbol_reg[3][3]  ( .D(n1283), .CK(clk), .RN(n1765), .Q(n2608), 
        .QN(n1574) );
  DFFRX1 \C1_symbol_reg[3][2]  ( .D(n1278), .CK(clk), .RN(n1761), .Q(n2609), 
        .QN(n1575) );
  DFFRX1 \C1_symbol_reg[3][1]  ( .D(n1273), .CK(clk), .RN(n1767), .Q(n2610), 
        .QN(n1571) );
  DFFRX1 \C1_symbol_reg[3][0]  ( .D(n1268), .CK(clk), .RN(n1759), .Q(n2611), 
        .QN(n1572) );
  DFFRX1 \C3_reg[2][5]  ( .D(n1213), .CK(clk), .RN(n1747), .Q(\C3[2][5] ), 
        .QN(n896) );
  DFFRX1 \C3_reg[2][1]  ( .D(n1225), .CK(clk), .RN(n1748), .Q(\C3[2][1] ), 
        .QN(n908) );
  DFFRX1 \C3_reg[2][4]  ( .D(n1216), .CK(clk), .RN(n1747), .Q(\C3[2][4] ), 
        .QN(n899) );
  DFFRX1 \C3_reg[1][6]  ( .D(n1209), .CK(clk), .RN(n1747), .Q(\C3[1][6] ), 
        .QN(n892) );
  DFFRX1 \C2_reg[3][3]  ( .D(n1242), .CK(clk), .RN(n1749), .Q(\C2[3][3] ), 
        .QN(n925) );
  DFFRX1 \C2_reg[3][6]  ( .D(n1254), .CK(clk), .RN(n1744), .Q(\C2[3][6] ), 
        .QN(n937) );
  DFFRX1 \C3_reg[0][1]  ( .D(n1223), .CK(clk), .RN(n1748), .QN(n906) );
  DFFRX1 \C1_reg[3][7]  ( .D(n1331), .CK(clk), .RN(n1762), .Q(\C1[3][7] ), 
        .QN(n1013) );
  DFFRX1 \C3_reg[0][5]  ( .D(n1211), .CK(clk), .RN(n1747), .QN(n894) );
  DFFRX1 \C3_reg[2][3]  ( .D(n1219), .CK(clk), .RN(n1747), .Q(\C3[2][3] ), 
        .QN(n902) );
  DFFRX1 \C1_reg[0][5]  ( .D(n1317), .CK(clk), .RN(n1762), .QN(n998) );
  DFFRX1 \C2_reg[0][5]  ( .D(n1251), .CK(clk), .RN(n1759), .QN(n931) );
  DFFRX1 \C2_reg[2][2]  ( .D(n1241), .CK(clk), .RN(n1749), .Q(\C2[2][2] ), 
        .QN(n922) );
  DFFRX1 \C3_reg[0][4]  ( .D(n1214), .CK(clk), .RN(n1747), .QN(n897) );
  DFFRX1 \C2_reg[2][3]  ( .D(n1245), .CK(clk), .RN(n1750), .Q(\C2[2][3] ), 
        .QN(n926) );
  DFFRX1 \symbol_value_reg[1][7]  ( .D(n1409), .CK(clk), .RN(n1761), .Q(
        \symbol_value[1][7] ), .QN(n1620) );
  DFFRX1 \C1_reg[1][7]  ( .D(n1329), .CK(clk), .RN(n1767), .Q(n1594), .QN(
        n1010) );
  DFFRX1 \C3_reg[1][2]  ( .D(n1221), .CK(clk), .RN(n1748), .Q(\C3[1][2] ), 
        .QN(n904) );
  DFFRX1 \C2_reg[1][4]  ( .D(n1248), .CK(clk), .RN(n1750), .Q(n1532), .QN(n928) );
  DFFRX1 \C2_reg[2][4]  ( .D(n1249), .CK(clk), .RN(n1750), .Q(\C2[2][4] ), 
        .QN(n930) );
  DFFRX1 \C2_reg[1][0]  ( .D(n1258), .CK(clk), .RN(n1757), .QN(n944) );
  DFFRX1 \symbol_value_reg[2][7]  ( .D(n1396), .CK(clk), .RN(n1759), .Q(
        \symbol_value[2][7] ), .QN(n1621) );
  DFFRX1 \C3_reg[1][3]  ( .D(n1218), .CK(clk), .RN(n1747), .Q(\C3[1][3] ), 
        .QN(n901) );
  DFFRX1 \C2_reg[1][2]  ( .D(n1240), .CK(clk), .RN(n1749), .Q(n1534), .QN(n920) );
  DFFRX2 \C2_reg[1][1]  ( .D(n1236), .CK(clk), .RN(n1749), .QN(n916) );
  DFFRX2 \symbol_value_reg[3][6]  ( .D(n1413), .CK(clk), .RN(n1761), .Q(
        \symbol_value[3][6] ), .QN(n1624) );
  DFFRX1 \C4_reg[0][2]  ( .D(n1201), .CK(clk), .RN(n1746), .Q(\C4[0][2] ), 
        .QN(n884) );
  DFFRX1 \C4_reg[0][4]  ( .D(n1197), .CK(clk), .RN(n1746), .Q(\C4[0][4] ), 
        .QN(n880) );
  DFFRX1 \C4_reg[1][2]  ( .D(n1200), .CK(clk), .RN(n1746), .Q(\C4[1][2] ), 
        .QN(n883) );
  DFFRX1 \C4_reg[1][4]  ( .D(n1196), .CK(clk), .RN(n1745), .Q(\C4[1][4] ), 
        .QN(n879) );
  DFFRX1 \C4_reg[0][5]  ( .D(n1195), .CK(clk), .RN(n1745), .Q(\C4[0][5] ), 
        .QN(n878) );
  DFFRX1 \C2_reg[3][2]  ( .D(n1238), .CK(clk), .RN(n1749), .Q(\C2[3][2] ), 
        .QN(n921) );
  DFFRX1 \C2_reg[2][0]  ( .D(n1263), .CK(clk), .RN(n1751), .Q(\C2[2][0] ), 
        .QN(n946) );
  DFFRX1 \C2_reg[2][1]  ( .D(n1237), .CK(clk), .RN(n1749), .Q(\C2[2][1] ), 
        .QN(n918) );
  DFFRX1 C4_sort_reg ( .D(n1422), .CK(clk), .RN(n1762), .Q(n2573), .QN(n1613)
         );
  DFFRX1 \C1_reg[2][6]  ( .D(n1324), .CK(clk), .RN(n1760), .Q(n1590), .QN(
        n1006) );
  DFFRX1 \C3_reg[1][5]  ( .D(n1212), .CK(clk), .RN(n1747), .Q(\C3[1][5] ), 
        .QN(n895) );
  DFFRX1 \C1_reg[2][7]  ( .D(n1330), .CK(clk), .RN(n1765), .Q(n1589), .QN(
        n1011) );
  DFFRX1 \C1_reg[2][2]  ( .D(n1304), .CK(clk), .RN(n1758), .Q(n1578), .QN(n986) );
  DFFRX1 \C1_reg[3][0]  ( .D(n1333), .CK(clk), .RN(n1752), .Q(\C1[3][0] ), 
        .QN(n1016) );
  DFFRX1 \C1_reg[2][4]  ( .D(n1314), .CK(clk), .RN(n1755), .Q(n1525), .QN(n996) );
  DFFRX1 \C1_reg[3][6]  ( .D(n1321), .CK(clk), .RN(n1759), .Q(\C1[3][6] ), 
        .QN(n1005) );
  DFFRX1 \C1_reg[2][3]  ( .D(n1309), .CK(clk), .RN(n1761), .Q(n1524), .QN(n991) );
  DFFRX1 \C1_reg[3][2]  ( .D(n1301), .CK(clk), .RN(n1764), .Q(\C1[3][2] ), 
        .QN(n985) );
  DFFRX1 \C1_reg[3][5]  ( .D(n1316), .CK(clk), .RN(n1759), .Q(\C1[3][5] ), 
        .QN(n1000) );
  DFFRX1 \C2_reg[2][5]  ( .D(n1253), .CK(clk), .RN(n1758), .Q(\C2[2][5] ), 
        .QN(n934) );
  DFFRX1 \C1_reg[3][1]  ( .D(n1296), .CK(clk), .RN(n1753), .Q(\C1[3][1] ), 
        .QN(n980) );
  DFFRX1 \symbol_value_reg[0][6]  ( .D(n1410), .CK(clk), .RN(n1767), .Q(
        \symbol_value[0][6] ), .QN(n1542) );
  DFFRX1 \C1_reg[3][3]  ( .D(n1306), .CK(clk), .RN(n1766), .Q(\C1[3][3] ), 
        .QN(n990) );
  DFFRX1 \C1_reg[3][4]  ( .D(n1311), .CK(clk), .RN(n1765), .Q(\C1[3][4] ), 
        .QN(n995) );
  DFFRX1 \C2_reg[1][5]  ( .D(n1252), .CK(clk), .RN(n1757), .Q(n1585), .QN(n932) );
  DFFRX1 \C1_reg[1][4]  ( .D(n1313), .CK(clk), .RN(n1763), .Q(n1526), .QN(n994) );
  DFFRX1 \C1_reg[1][0]  ( .D(n1327), .CK(clk), .RN(n1764), .QN(n1008) );
  DFFRX1 \symbol_value_reg[0][7]  ( .D(n1408), .CK(clk), .RN(n1762), .Q(
        \symbol_value[0][7] ), .QN(n1610) );
  DFFRX1 \C1_reg[1][6]  ( .D(n1323), .CK(clk), .RN(n1766), .Q(n1582), .QN(
        n1004) );
  DFFRX1 \symbol_value_reg[0][3]  ( .D(n1338), .CK(clk), .RN(n1751), .Q(
        \symbol_value[0][3] ), .QN(n1616) );
  DFFRX1 \symbol_value_reg[0][4]  ( .D(n1334), .CK(clk), .RN(n1741), .Q(
        \symbol_value[0][4] ), .QN(n1615) );
  DFFRX1 \C1_reg[1][2]  ( .D(n1303), .CK(clk), .RN(n1767), .Q(n1533), .QN(n984) );
  DFFRX2 \sort_stage_reg[2]  ( .D(n1428), .CK(clk), .RN(n1767), .Q(
        sort_stage[2]) );
  DFFRX2 \C1_reg[1][1]  ( .D(n1298), .CK(clk), .RN(n1763), .QN(n979) );
  DFFRX2 \symbol_value_reg[4][7]  ( .D(n1417), .CK(clk), .RN(n1762), .Q(
        \symbol_value[4][7] ), .QN(n1609) );
  DFFRX2 \symbol_value_reg[1][6]  ( .D(n1411), .CK(clk), .RN(n1765), .Q(
        \symbol_value[1][6] ), .QN(n1652) );
  DFFRX2 \sort_stage_reg[0]  ( .D(n1420), .CK(clk), .RN(n1758), .Q(
        sort_stage[0]), .QN(n1688) );
  DFFRX1 \C1_reg[2][0]  ( .D(n1325), .CK(clk), .RN(n1756), .Q(n1579), .QN(
        n1014) );
  DFFRX1 \C1_reg[2][1]  ( .D(n1299), .CK(clk), .RN(n1766), .Q(n1523), .QN(n981) );
  DFFRX1 \symbol_value_reg[0][0]  ( .D(n1343), .CK(clk), .RN(n1742), .Q(
        \symbol_value[0][0] ), .QN(n1596) );
  DFFRX1 \C1_reg[2][5]  ( .D(n1319), .CK(clk), .RN(n1762), .Q(n1577), .QN(
        n1001) );
  DFFRX1 \sort_stage_reg[1]  ( .D(n1419), .CK(clk), .RN(n1760), .Q(
        sort_stage[1]), .QN(n1581) );
  DFFRX1 \symbol_value_reg[0][1]  ( .D(n1348), .CK(clk), .RN(n1754), .Q(
        \symbol_value[0][1] ), .QN(n1535) );
  DFFRX1 \symbol_value_reg[1][2]  ( .D(n1353), .CK(clk), .RN(n1751), .Q(
        \symbol_value[1][2] ), .QN(n1527) );
  DFFRX1 \C1_reg[1][5]  ( .D(n1318), .CK(clk), .RN(n1760), .Q(n1584), .QN(n999) );
  DFFRX1 \symbol_value_reg[1][4]  ( .D(n1397), .CK(clk), .RN(n1764), .Q(
        \symbol_value[1][4] ), .QN(n1539) );
  DFFRX1 \symbol_value_reg[0][5]  ( .D(n1407), .CK(clk), .RN(n1754), .Q(
        \symbol_value[0][5] ), .QN(n1597) );
  DFFRX2 \symbol_value_reg[1][1]  ( .D(n1349), .CK(clk), .RN(n1747), .Q(
        \symbol_value[1][1] ), .QN(n1653) );
  DFFRX2 \symbol_value_reg[4][2]  ( .D(n1356), .CK(clk), .RN(n1760), .Q(
        \symbol_value[4][2] ), .QN(n1685) );
  DFFRX1 \symbol_reg[5][0]  ( .D(n1392), .CK(clk), .RN(n1766), .Q(
        \symbol[5][0] ), .QN(n1655) );
  DFFRX1 \symbol_reg[5][1]  ( .D(n1386), .CK(clk), .RN(n1760), .Q(
        \symbol[5][1] ), .QN(n1656) );
  DFFRX1 \symbol_reg[5][2]  ( .D(n1380), .CK(clk), .RN(n1758), .Q(
        \symbol[5][2] ), .QN(n1657) );
  DFFRX1 \symbol_reg[5][3]  ( .D(n1374), .CK(clk), .RN(n1762), .Q(
        \symbol[5][3] ), .QN(n1658) );
  DFFRX1 \symbol_reg[5][4]  ( .D(n1368), .CK(clk), .RN(n1760), .Q(
        \symbol[5][4] ), .QN(n1659) );
  DFFRX1 \symbol_reg[4][0]  ( .D(n1393), .CK(clk), .RN(n1757), .Q(
        \symbol[4][0] ), .QN(n1493) );
  DFFRX1 \symbol_reg[4][1]  ( .D(n1387), .CK(clk), .RN(n1758), .Q(
        \symbol[4][1] ), .QN(n1494) );
  DFFRX1 \symbol_reg[4][2]  ( .D(n1381), .CK(clk), .RN(n1764), .Q(
        \symbol[4][2] ), .QN(n1495) );
  DFFRX1 \symbol_reg[4][3]  ( .D(n1375), .CK(clk), .RN(n1761), .Q(
        \symbol[4][3] ), .QN(n1521) );
  DFFSX1 \symbol_reg[4][4]  ( .D(n1369), .CK(clk), .SN(n1756), .Q(
        \symbol[4][4] ), .QN(n1496) );
  DFFRX1 \state_reg[2]  ( .D(n1423), .CK(clk), .RN(n1757), .Q(state[2]), .QN(
        n1586) );
  DFFRX1 \state_reg[0]  ( .D(n1427), .CK(clk), .RN(n1760), .Q(state[0]), .QN(
        n1580) );
  DFFRX1 \symbol_value_reg[5][7]  ( .D(n1416), .CK(clk), .RN(n1756), .Q(
        \symbol_value[5][7] ), .QN(n1623) );
  DFFRX1 \symbol_value_reg[2][0]  ( .D(n1345), .CK(clk), .RN(n1741), .Q(
        \symbol_value[2][0] ), .QN(n1606) );
  DFFRX1 \symbol_value_reg[2][3]  ( .D(n1351), .CK(clk), .RN(n1742), .Q(
        \symbol_value[2][3] ), .QN(n1538) );
  DFFRX1 \symbol_value_reg[2][4]  ( .D(n1398), .CK(clk), .RN(n1760), .Q(
        \symbol_value[2][4] ), .QN(n1541) );
  DFFRX1 \symbol_value_reg[2][2]  ( .D(n1354), .CK(clk), .RN(n1756), .Q(
        \symbol_value[2][2] ), .QN(n1605) );
  DFFRX1 \symbol_value_reg[1][5]  ( .D(n1406), .CK(clk), .RN(n2619), .Q(
        \symbol_value[1][5] ), .QN(n1604) );
  DFFRX1 \symbol_value_reg[2][5]  ( .D(n1405), .CK(clk), .RN(n2619), .Q(
        \symbol_value[2][5] ), .QN(n1592) );
  DFFRX1 \symbol_value_reg[2][1]  ( .D(n1350), .CK(clk), .RN(n1746), .Q(
        \symbol_value[2][1] ), .QN(n1531) );
  DFFRX1 \symbol_value_reg[5][0]  ( .D(n1341), .CK(clk), .RN(n1746), .Q(
        \symbol_value[5][0] ) );
  DFFRX1 \symbol_value_reg[3][3]  ( .D(n1358), .CK(clk), .RN(n1756), .Q(
        \symbol_value[3][3] ), .QN(n1540) );
  DFFRX1 \symbol_value_reg[4][6]  ( .D(n1414), .CK(clk), .RN(n1759), .Q(
        \symbol_value[4][6] ), .QN(n1529) );
  DFFRX1 \symbol_value_reg[4][3]  ( .D(n1357), .CK(clk), .RN(n1745), .Q(
        \symbol_value[4][3] ), .QN(n1591) );
  DFFRX1 \symbol_value_reg[4][4]  ( .D(n1400), .CK(clk), .RN(n1758), .Q(
        \symbol_value[4][4] ), .QN(n1593) );
  DFFRX1 \symbol_value_reg[5][6]  ( .D(n1415), .CK(clk), .RN(n1763), .Q(
        \symbol_value[5][6] ) );
  DFFRX1 \symbol_value_reg[5][4]  ( .D(n1401), .CK(clk), .RN(n1767), .Q(
        \symbol_value[5][4] ) );
  DFFRX1 \symbol_value_reg[4][1]  ( .D(n1340), .CK(clk), .RN(n1745), .Q(
        \symbol_value[4][1] ), .QN(n1528) );
  DFFRX1 \symbol_value_reg[1][3]  ( .D(n1352), .CK(clk), .RN(n1743), .Q(
        \symbol_value[1][3] ), .QN(n1588) );
  DFFRX1 \symbol_value_reg[0][2]  ( .D(n1337), .CK(clk), .RN(n1743), .Q(
        \symbol_value[0][2] ), .QN(n1639) );
  DFFRX1 \symbol_value_reg[4][5]  ( .D(n1403), .CK(clk), .RN(n1759), .Q(
        \symbol_value[4][5] ), .QN(n1530) );
  DFFRX1 \symbol_value_reg[5][2]  ( .D(n1336), .CK(clk), .RN(n1744), .Q(
        \symbol_value[5][2] ), .QN(n1545) );
  DFFRX1 \symbol_value_reg[5][5]  ( .D(n1402), .CK(clk), .RN(n1761), .Q(
        \symbol_value[5][5] ) );
  DFFRX1 \symbol_value_reg[5][1]  ( .D(n1339), .CK(clk), .RN(n1755), .Q(
        \symbol_value[5][1] ) );
  DFFRX1 C3_sort_reg ( .D(n1421), .CK(clk), .RN(n1765), .Q(n2586), .QN(n1587)
         );
  DFFRX1 \state_reg[1]  ( .D(n1425), .CK(clk), .RN(n1749), .Q(state[1]), .QN(
        n1583) );
  DFFRX2 C1_sort_reg ( .D(n1426), .CK(clk), .RN(n1765), .Q(n2618), .QN(n1626)
         );
  DFFRX2 C2_sort_reg ( .D(n1429), .CK(clk), .RN(n1747), .Q(n2599), .QN(n1614)
         );
  DFFRX1 \symbol_value_reg[1][0]  ( .D(n1344), .CK(clk), .RN(n1754), .Q(
        \symbol_value[1][0] ), .QN(n1654) );
  DFFRX1 \symbol_value_reg[3][7]  ( .D(n1395), .CK(clk), .RN(n1744), .Q(
        \symbol_value[3][7] ), .QN(n1625) );
  DFFRX1 \symbol_value_reg[2][6]  ( .D(n1412), .CK(clk), .RN(n1762), .Q(
        \symbol_value[2][6] ), .QN(n1622) );
  DFFRX1 \symbol_value_reg[5][3]  ( .D(n1335), .CK(clk), .RN(n1753), .Q(
        \symbol_value[5][3] ), .QN(n1619) );
  DFFRX1 \symbol_value_reg[3][0]  ( .D(n1346), .CK(clk), .RN(n1744), .Q(
        \symbol_value[3][0] ), .QN(n1618) );
  DFFRX1 \C2_reg[1][6]  ( .D(n1256), .CK(clk), .RN(n1757), .Q(n1617), .QN(n936) );
  DFFRX1 \symbol_value_reg[3][2]  ( .D(n1355), .CK(clk), .RN(n1750), .Q(
        \symbol_value[3][2] ), .QN(n1612) );
  DFFRX1 \symbol_value_reg[3][4]  ( .D(n1399), .CK(clk), .RN(n1759), .Q(
        \symbol_value[3][4] ), .QN(n1611) );
  DFFRX1 \symbol_value_reg[4][0]  ( .D(n1342), .CK(clk), .RN(n1757), .Q(
        \symbol_value[4][0] ), .QN(n1608) );
  DFFRX1 \C2_reg[1][3]  ( .D(n1244), .CK(clk), .RN(n1749), .Q(n1601), .QN(n924) );
  DFFRX1 \C1_reg[1][3]  ( .D(n1308), .CK(clk), .RN(n1748), .Q(n1600), .QN(n989) );
  DFFRX1 \symbol_value_reg[3][1]  ( .D(n1347), .CK(clk), .RN(n1748), .Q(
        \symbol_value[3][1] ), .QN(n1544) );
  DFFRX1 \symbol_value_reg[3][5]  ( .D(n1404), .CK(clk), .RN(n1760), .Q(
        \symbol_value[3][5] ), .QN(n1543) );
  NOR2X2 U1152 ( .A(n1830), .B(gray_valid), .Y(n1478) );
  NAND2X1 U1153 ( .A(n2573), .B(n1739), .Y(n1480) );
  NAND2X1 U1154 ( .A(n1613), .B(n1739), .Y(n1481) );
  OAI21X1 U1155 ( .A0(n2276), .A1(n1632), .B0(n1709), .Y(n2272) );
  OAI21X1 U1156 ( .A0(n2276), .A1(n2524), .B0(n1709), .Y(n2283) );
  OAI21X1 U1157 ( .A0(n2309), .A1(n1633), .B0(n1710), .Y(n2305) );
  OAI21X1 U1158 ( .A0(n2309), .A1(n2533), .B0(n1710), .Y(n2316) );
  OAI21X1 U1159 ( .A0(n2342), .A1(n1634), .B0(n1711), .Y(n2338) );
  OAI21X2 U1160 ( .A0(\symbol[5][4] ), .A1(\symbol[4][4] ), .B0(n2253), .Y(
        n2271) );
  OAI21X1 U1161 ( .A0(n2342), .A1(n2542), .B0(n1711), .Y(n2349) );
  OAI21X1 U1162 ( .A0(n2375), .A1(n1635), .B0(n1712), .Y(n2371) );
  OAI21X1 U1163 ( .A0(n2487), .A1(n2560), .B0(n1727), .Y(n2483) );
  AND2X2 U1164 ( .A(n1693), .B(n1891), .Y(n1855) );
  OAI211X4 U1165 ( .A0(n1975), .A1(n1976), .B0(n1830), .C0(n1834), .Y(n1891)
         );
  OAI21X2 U1166 ( .A0(\symbol[5][3] ), .A1(\symbol[4][3] ), .B0(n2253), .Y(
        n2304) );
  OA21X2 U1167 ( .A0(n1708), .A1(n1637), .B0(n1707), .Y(n2233) );
  NAND2X2 U1168 ( .A(n1824), .B(n1614), .Y(n2258) );
  NOR3X2 U1169 ( .A(sort_stage[1]), .B(sort_stage[2]), .C(n1830), .Y(n1843) );
  OAI21X1 U1170 ( .A0(n2375), .A1(n2551), .B0(n1712), .Y(n2382) );
  OAI21X1 U1171 ( .A0(n2487), .A1(n1636), .B0(n1727), .Y(n2493) );
  NOR2X2 U1172 ( .A(gray_valid), .B(n1867), .Y(n1868) );
  NOR2X2 U1173 ( .A(n1768), .B(n1855), .Y(n1857) );
  OAI21X2 U1174 ( .A0(\symbol[5][2] ), .A1(\symbol[4][2] ), .B0(n2253), .Y(
        n2337) );
  OA21X2 U1175 ( .A0(n1708), .A1(n2515), .B0(n1707), .Y(n2244) );
  NAND2X2 U1176 ( .A(n1844), .B(n1587), .Y(n2257) );
  CLKINVX2 U1177 ( .A(n2184), .Y(n2153) );
  NAND2X2 U1178 ( .A(n2504), .B(n1580), .Y(n1828) );
  AND2X2 U1179 ( .A(n1694), .B(n1898), .Y(n1867) );
  OAI211X4 U1180 ( .A0(n1992), .A1(n1993), .B0(n1830), .C0(n1834), .Y(n1898)
         );
  NOR2X2 U1181 ( .A(gray_valid), .B(n1855), .Y(n1856) );
  NOR2X2 U1182 ( .A(n1768), .B(n1867), .Y(n1869) );
  NOR2BX2 U1183 ( .AN(n1689), .B(n1887), .Y(n1861) );
  NOR2BX2 U1184 ( .AN(n1690), .B(n1894), .Y(n1863) );
  NOR2BX2 U1185 ( .AN(n1691), .B(n1897), .Y(n1865) );
  NOR2BX2 U1186 ( .AN(n1692), .B(n1890), .Y(n1852) );
  OAI21X2 U1187 ( .A0(\symbol[5][1] ), .A1(\symbol[4][1] ), .B0(n2253), .Y(
        n2370) );
  OAI21X2 U1188 ( .A0(\symbol[5][0] ), .A1(\symbol[4][0] ), .B0(n2253), .Y(
        n2482) );
  NOR2X2 U1189 ( .A(n1822), .B(n2618), .Y(n2253) );
  INVX1 U1190 ( .A(n1828), .Y(n1846) );
  INVX1 U1191 ( .A(n2482), .Y(n2487) );
  INVX1 U1192 ( .A(n2370), .Y(n2375) );
  INVX1 U1193 ( .A(n2337), .Y(n2342) );
  INVX1 U1194 ( .A(n2304), .Y(n2309) );
  INVX1 U1195 ( .A(n2271), .Y(n2276) );
  INVX1 U1196 ( .A(n1843), .Y(n1847) );
  INVX1 U1197 ( .A(n2253), .Y(n2084) );
  NAND2XL U1198 ( .A(n1626), .B(n1706), .Y(n2062) );
  MXI2XL U1199 ( .A(n1496), .B(n1659), .S0(n1891), .Y(n1368) );
  MXI2XL U1200 ( .A(n1521), .B(n1658), .S0(n1891), .Y(n1374) );
  MXI2XL U1201 ( .A(n1495), .B(n1657), .S0(n1891), .Y(n1380) );
  MXI2XL U1202 ( .A(n1494), .B(n1656), .S0(n1891), .Y(n1386) );
  MXI2XL U1203 ( .A(n1493), .B(n1655), .S0(n1891), .Y(n1392) );
  MXI2XL U1204 ( .A(n1564), .B(n1684), .S0(n1891), .Y(n1362) );
  MXI2XL U1205 ( .A(n1487), .B(n1646), .S0(n1898), .Y(n1359) );
  MXI2XL U1206 ( .A(n1516), .B(n1647), .S0(n1898), .Y(n1365) );
  MXI2XL U1207 ( .A(n1517), .B(n1648), .S0(n1898), .Y(n1371) );
  MXI2XL U1208 ( .A(n1518), .B(n1649), .S0(n1898), .Y(n1377) );
  MXI2XL U1209 ( .A(n1519), .B(n1650), .S0(n1898), .Y(n1383) );
  MXI2XL U1210 ( .A(n1520), .B(n1651), .S0(n1898), .Y(n1389) );
  NAND2XL U1211 ( .A(n1626), .B(n1822), .Y(n1426) );
  NAND2XL U1212 ( .A(n1614), .B(n1728), .Y(n1429) );
  NAND2XL U1213 ( .A(n1613), .B(n1828), .Y(n1422) );
  AOI21XL U1214 ( .A0(n2482), .A1(n2478), .B0(n2493), .Y(n2492) );
  AOI21XL U1215 ( .A0(n2482), .A1(n2478), .B0(n2483), .Y(n2481) );
  AOI21XL U1216 ( .A0(n2370), .A1(n2367), .B0(n2382), .Y(n2381) );
  AOI21XL U1217 ( .A0(n2370), .A1(n2367), .B0(n2371), .Y(n2369) );
  AOI21XL U1218 ( .A0(n2337), .A1(n2334), .B0(n2349), .Y(n2348) );
  AOI21XL U1219 ( .A0(n2337), .A1(n2334), .B0(n2338), .Y(n2336) );
  AOI21XL U1220 ( .A0(n2304), .A1(n2301), .B0(n2316), .Y(n2315) );
  AOI21XL U1221 ( .A0(n2304), .A1(n2301), .B0(n2305), .Y(n2303) );
  AOI21XL U1222 ( .A0(n2271), .A1(n2268), .B0(n2283), .Y(n2282) );
  AOI21XL U1223 ( .A0(n2271), .A1(n2268), .B0(n2272), .Y(n2270) );
  AOI21XL U1224 ( .A0(n1784), .A1(n2482), .B0(n2493), .Y(n2494) );
  AOI21XL U1225 ( .A0(n1784), .A1(n2482), .B0(n2483), .Y(n2484) );
  AOI21XL U1226 ( .A0(n1788), .A1(n2370), .B0(n2382), .Y(n2383) );
  AOI21XL U1227 ( .A0(n1788), .A1(n2370), .B0(n2371), .Y(n2372) );
  AOI21XL U1228 ( .A0(n1792), .A1(n2337), .B0(n2349), .Y(n2350) );
  AOI21XL U1229 ( .A0(n1792), .A1(n2337), .B0(n2338), .Y(n2339) );
  AOI21XL U1230 ( .A0(n1796), .A1(n2304), .B0(n2316), .Y(n2317) );
  AOI21XL U1231 ( .A0(n1796), .A1(n2304), .B0(n2305), .Y(n2306) );
  AOI21XL U1232 ( .A0(n1800), .A1(n2271), .B0(n2283), .Y(n2284) );
  AOI21XL U1233 ( .A0(n1800), .A1(n2271), .B0(n2272), .Y(n2273) );
  AOI2BB1XL U1234 ( .A0N(n1785), .A1N(n2487), .B0(n2493), .Y(n2495) );
  AOI2BB1XL U1235 ( .A0N(n1785), .A1N(n2487), .B0(n2483), .Y(n2486) );
  AOI2BB1XL U1236 ( .A0N(n1789), .A1N(n2375), .B0(n2382), .Y(n2384) );
  AOI2BB1XL U1237 ( .A0N(n1789), .A1N(n2375), .B0(n2371), .Y(n2374) );
  AOI2BB1XL U1238 ( .A0N(n1793), .A1N(n2342), .B0(n2349), .Y(n2351) );
  AOI2BB1XL U1239 ( .A0N(n1793), .A1N(n2342), .B0(n2338), .Y(n2341) );
  AOI2BB1XL U1240 ( .A0N(n1797), .A1N(n2309), .B0(n2316), .Y(n2318) );
  AOI2BB1XL U1241 ( .A0N(n1797), .A1N(n2309), .B0(n2305), .Y(n2308) );
  AOI2BB1XL U1242 ( .A0N(n1801), .A1N(n2276), .B0(n2283), .Y(n2285) );
  AOI2BB1XL U1243 ( .A0N(n1801), .A1N(n2276), .B0(n2272), .Y(n2275) );
  OAI211XL U1244 ( .A0(\symbol[4][0] ), .A1(n2482), .B0(n2496), .C0(n2497), 
        .Y(n1024) );
  OAI211XL U1245 ( .A0(\symbol[4][1] ), .A1(n2370), .B0(n2376), .C0(n2377), 
        .Y(n1064) );
  OAI211XL U1246 ( .A0(\symbol[4][2] ), .A1(n2337), .B0(n2343), .C0(n2344), 
        .Y(n1092) );
  OAI211XL U1247 ( .A0(\symbol[4][3] ), .A1(n2304), .B0(n2310), .C0(n2311), 
        .Y(n1120) );
  OAI211XL U1248 ( .A0(\symbol[4][4] ), .A1(n2271), .B0(n2277), .C0(n2278), 
        .Y(n1148) );
  OA22XL U1249 ( .A0(n2257), .A1(n2440), .B0(n2258), .B1(n2392), .Y(n2502) );
  OA22XL U1250 ( .A0(n2257), .A1(n2362), .B0(n2258), .B1(n2359), .Y(n2391) );
  OAI211XL U1251 ( .A0(n2331), .A1(n2254), .B0(n2357), .C0(n2358), .Y(n2354)
         );
  OA22XL U1252 ( .A0(n2257), .A1(n2329), .B0(n2258), .B1(n2326), .Y(n2358) );
  OAI211XL U1253 ( .A0(n2298), .A1(n2254), .B0(n2324), .C0(n2325), .Y(n2321)
         );
  OA22XL U1254 ( .A0(n2257), .A1(n2296), .B0(n2258), .B1(n2293), .Y(n2325) );
  OAI211XL U1255 ( .A0(n2265), .A1(n2254), .B0(n2291), .C0(n2292), .Y(n2288)
         );
  OA22XL U1256 ( .A0(n2257), .A1(n2263), .B0(n2258), .B1(n2260), .Y(n2292) );
  NAND2XL U1257 ( .A(n1843), .B(n2086), .Y(n2081) );
  AOI22XL U1258 ( .A0(n2010), .A1(n1523), .B0(n2011), .B1(\symbol_value[3][1] ), .Y(n2054) );
  AOI22XL U1259 ( .A0(n2609), .A1(n1696), .B0(n2615), .B1(n2059), .Y(n2072) );
  AOI22XL U1260 ( .A0(n2608), .A1(n1696), .B0(n2614), .B1(n2059), .Y(n2068) );
  AOI22XL U1261 ( .A0(n2607), .A1(n1696), .B0(n2613), .B1(n2059), .Y(n2064) );
  AOI22XL U1262 ( .A0(n2606), .A1(n1696), .B0(n2612), .B1(n2059), .Y(n2058) );
  MXI2XL U1263 ( .A(n1953), .B(n1528), .S0(n1852), .Y(n1340) );
  MXI2XL U1264 ( .A(n1900), .B(n1591), .S0(n1852), .Y(n1357) );
  MXI2XL U1265 ( .A(n1879), .B(n1593), .S0(n1852), .Y(n1400) );
  MXI2XL U1266 ( .A(n1876), .B(n1530), .S0(n1852), .Y(n1403) );
  MXI2XL U1267 ( .A(n1859), .B(n1529), .S0(n1852), .Y(n1414) );
  OAI211XL U1268 ( .A0(n2225), .A1(n2254), .B0(n2255), .C0(n2256), .Y(n2249)
         );
  OA22XL U1269 ( .A0(n2257), .A1(n2223), .B0(n2258), .B1(n2220), .Y(n2256) );
  AOI2BB2XL U1270 ( .B0(N1726), .B1(n2153), .A0N(n2154), .A1N(n946), .Y(n2152)
         );
  AOI2BB2XL U1271 ( .B0(N1733), .B1(n2153), .A0N(n2154), .A1N(n943), .Y(n2183)
         );
  AOI2BB2XL U1272 ( .B0(N1727), .B1(n2153), .A0N(n2154), .A1N(n918), .Y(n2182)
         );
  AOI2BB2XL U1273 ( .B0(N1728), .B1(n2153), .A0N(n2154), .A1N(n922), .Y(n2179)
         );
  AOI2BB2XL U1274 ( .B0(N1729), .B1(n2153), .A0N(n2154), .A1N(n926), .Y(n2176)
         );
  AOI2BB2XL U1275 ( .B0(N1730), .B1(n2153), .A0N(n2154), .A1N(n930), .Y(n2173)
         );
  AOI2BB2XL U1276 ( .B0(N1731), .B1(n2153), .A0N(n2154), .A1N(n934), .Y(n2170)
         );
  AOI2BB2XL U1277 ( .B0(N1732), .B1(n2153), .A0N(n2154), .A1N(n938), .Y(n2167)
         );
  OAI2BB1XL U1278 ( .A0N(\symbol_value[4][0] ), .A1N(n1856), .B0(n1952), .Y(
        n1341) );
  MXI2XL U1279 ( .A(n1857), .B(n1855), .S0(\symbol_value[5][0] ), .Y(n1952) );
  OAI2BB1XL U1280 ( .A0N(\symbol_value[1][0] ), .A1N(n1868), .B0(n1950), .Y(
        n1343) );
  MXI2XL U1281 ( .A(n1867), .B(n1869), .S0(n1596), .Y(n1950) );
  AOI211XL U1282 ( .A0(n980), .A1(n1523), .B0(n1579), .C0(n1016), .Y(n2098) );
  NOR2XL U1283 ( .A(n980), .B(n1523), .Y(n2099) );
  AND2XL U1284 ( .A(n979), .B(n1523), .Y(n2115) );
  OAI211XL U1285 ( .A0(n1523), .A1(n979), .B0(n1008), .C0(n1579), .Y(n2116) );
  AND2XL U1286 ( .A(n2254), .B(n2475), .Y(n1686) );
  AOI33XL U1287 ( .A0(n1843), .A1(n1844), .A2(n2586), .B0(n1845), .B1(n1846), 
        .B2(n2573), .Y(n1839) );
  MXI2XL U1288 ( .A(n1901), .B(n1685), .S0(n1852), .Y(n1356) );
  MXI2XL U1289 ( .A(n1884), .B(n1625), .S0(n1861), .Y(n1395) );
  MXI2XL U1290 ( .A(n1851), .B(n1609), .S0(n1852), .Y(n1417) );
  MXI2XL U1291 ( .A(n1910), .B(n1544), .S0(n1861), .Y(n1347) );
  MXI2XL U1292 ( .A(n1908), .B(n1653), .S0(n1865), .Y(n1349) );
  MXI2XL U1293 ( .A(n1902), .B(n1612), .S0(n1861), .Y(n1355) );
  MXI2XL U1294 ( .A(n1880), .B(n1611), .S0(n1861), .Y(n1399) );
  MXI2XL U1295 ( .A(n1875), .B(n1543), .S0(n1861), .Y(n1404) );
  MXI2XL U1296 ( .A(n1864), .B(n1652), .S0(n1865), .Y(n1411) );
  MXI2XL U1297 ( .A(n1862), .B(n1622), .S0(n1863), .Y(n1412) );
  MXI2XL U1298 ( .A(n1860), .B(n1624), .S0(n1861), .Y(n1413) );
  MXI2XL U1299 ( .A(n1883), .B(n1621), .S0(n1863), .Y(n1396) );
  MXI2XL U1300 ( .A(n1870), .B(n1620), .S0(n1865), .Y(n1409) );
  MXI2XL U1301 ( .A(n1907), .B(n1531), .S0(n1863), .Y(n1350) );
  MXI2XL U1302 ( .A(n1906), .B(n1538), .S0(n1863), .Y(n1351) );
  MXI2XL U1303 ( .A(n1905), .B(n1588), .S0(n1865), .Y(n1352) );
  MXI2XL U1304 ( .A(n1904), .B(n1527), .S0(n1865), .Y(n1353) );
  MXI2XL U1305 ( .A(n1903), .B(n1605), .S0(n1863), .Y(n1354) );
  MXI2XL U1306 ( .A(n1899), .B(n1540), .S0(n1861), .Y(n1358) );
  MXI2XL U1307 ( .A(n1882), .B(n1539), .S0(n1865), .Y(n1397) );
  MXI2XL U1308 ( .A(n1881), .B(n1541), .S0(n1863), .Y(n1398) );
  MXI2XL U1309 ( .A(n1874), .B(n1592), .S0(n1863), .Y(n1405) );
  MXI2XL U1310 ( .A(n1873), .B(n1604), .S0(n1865), .Y(n1406) );
  NAND2XL U1311 ( .A(n1843), .B(n2411), .Y(n2394) );
  NOR3XL U1312 ( .A(n1626), .B(sort_stage[2]), .C(n1822), .Y(n1835) );
  AOI211XL U1313 ( .A0(n1838), .A1(n1847), .B0(n1614), .C0(n1728), .Y(n1836)
         );
  CLKINVX1 U1314 ( .A(gray_valid), .Y(n1768) );
  CLKBUFX3 U1315 ( .A(n1759), .Y(n1751) );
  CLKBUFX3 U1316 ( .A(n1759), .Y(n1752) );
  CLKBUFX3 U1317 ( .A(n1756), .Y(n1753) );
  CLKBUFX3 U1318 ( .A(n1758), .Y(n1754) );
  CLKBUFX3 U1319 ( .A(n1758), .Y(n1755) );
  CLKBUFX3 U1320 ( .A(n1761), .Y(n1747) );
  CLKBUFX3 U1321 ( .A(n1761), .Y(n1748) );
  CLKBUFX3 U1322 ( .A(n1760), .Y(n1749) );
  CLKBUFX3 U1323 ( .A(n1760), .Y(n1750) );
  CLKBUFX3 U1324 ( .A(n1763), .Y(n1742) );
  CLKBUFX3 U1325 ( .A(n1764), .Y(n1743) );
  CLKBUFX3 U1326 ( .A(n1766), .Y(n1744) );
  CLKBUFX3 U1327 ( .A(n1762), .Y(n1745) );
  CLKBUFX3 U1328 ( .A(n1762), .Y(n1746) );
  CLKBUFX3 U1329 ( .A(n1763), .Y(n1741) );
  CLKBUFX3 U1330 ( .A(n1766), .Y(n1756) );
  CLKBUFX3 U1331 ( .A(n1765), .Y(n1759) );
  CLKBUFX3 U1332 ( .A(n1745), .Y(n1758) );
  CLKBUFX3 U1333 ( .A(n1765), .Y(n1761) );
  CLKBUFX3 U1334 ( .A(n1765), .Y(n1760) );
  CLKBUFX3 U1335 ( .A(n1750), .Y(n1757) );
  CLKBUFX3 U1336 ( .A(n1481), .Y(n1735) );
  CLKBUFX3 U1337 ( .A(n1478), .Y(n1732) );
  CLKBUFX3 U1338 ( .A(n1764), .Y(n1762) );
  CLKBUFX3 U1339 ( .A(n1764), .Y(n1763) );
  CLKBUFX3 U1340 ( .A(n1767), .Y(n1765) );
  CLKBUFX3 U1341 ( .A(n1786), .Y(n1727) );
  CLKINVX1 U1342 ( .A(n2476), .Y(n1786) );
  CLKBUFX3 U1343 ( .A(n1790), .Y(n1712) );
  CLKINVX1 U1344 ( .A(n2365), .Y(n1790) );
  CLKBUFX3 U1345 ( .A(n1794), .Y(n1711) );
  CLKINVX1 U1346 ( .A(n2332), .Y(n1794) );
  CLKBUFX3 U1347 ( .A(n1798), .Y(n1710) );
  CLKINVX1 U1348 ( .A(n2299), .Y(n1798) );
  CLKBUFX3 U1349 ( .A(n1802), .Y(n1709) );
  CLKINVX1 U1350 ( .A(n2266), .Y(n1802) );
  CLKBUFX3 U1351 ( .A(n1806), .Y(n1707) );
  CLKINVX1 U1352 ( .A(n2226), .Y(n1806) );
  CLKBUFX3 U1353 ( .A(n2014), .Y(n1705) );
  CLKINVX1 U1354 ( .A(n2062), .Y(n2014) );
  CLKBUFX3 U1355 ( .A(n1480), .Y(n1738) );
  CLKBUFX3 U1356 ( .A(n1739), .Y(n1740) );
  CLKBUFX3 U1357 ( .A(n1481), .Y(n1736) );
  CLKBUFX3 U1358 ( .A(n1853), .Y(n1734) );
  CLKBUFX3 U1359 ( .A(n1478), .Y(n1731) );
  CLKBUFX3 U1360 ( .A(n1766), .Y(n1764) );
  CLKBUFX3 U1361 ( .A(n1767), .Y(n1766) );
  CLKBUFX3 U1362 ( .A(n2020), .Y(n1696) );
  NOR3XL U1363 ( .A(n2059), .B(n2083), .C(n1626), .Y(n2020) );
  CLKBUFX3 U1364 ( .A(n2021), .Y(n1699) );
  NAND2X1 U1365 ( .A(n2084), .B(n2085), .Y(n2021) );
  CLKBUFX3 U1366 ( .A(n2231), .Y(n1708) );
  NOR2X1 U1367 ( .A(n2084), .B(n2061), .Y(n2231) );
  CLKBUFX3 U1368 ( .A(n2027), .Y(n1703) );
  NAND2XL U1369 ( .A(n1626), .B(n1704), .Y(n2027) );
  AND2X2 U1370 ( .A(n1918), .B(n1913), .Y(n1894) );
  AND2X2 U1371 ( .A(n1912), .B(n1913), .Y(n1887) );
  CLKAND2X3 U1372 ( .A(n1695), .B(n1626), .Y(n2011) );
  CLKAND2X3 U1373 ( .A(n1713), .B(n1614), .Y(n2149) );
  CLKBUFX3 U1374 ( .A(n2147), .Y(n1713) );
  AO21X1 U1375 ( .A0(n1824), .A1(n2395), .B0(n1714), .Y(n2147) );
  CLKBUFX3 U1376 ( .A(n2193), .Y(n1724) );
  NAND2BX1 U1377 ( .AN(n1726), .B(n2441), .Y(n2193) );
  CLKBUFX3 U1378 ( .A(n2008), .Y(n1695) );
  AO21X1 U1379 ( .A0(n1825), .A1(n2080), .B0(n1706), .Y(n2008) );
  CLKBUFX3 U1380 ( .A(n2185), .Y(n1721) );
  NAND2XL U1381 ( .A(n2257), .B(n2441), .Y(n2185) );
  CLKBUFX3 U1382 ( .A(n2160), .Y(n1717) );
  AO21X1 U1383 ( .A0(n1824), .A1(n2395), .B0(n1719), .Y(n2160) );
  CLKBUFX3 U1384 ( .A(n2026), .Y(n1702) );
  AO21X1 U1385 ( .A0(n1825), .A1(n2083), .B0(n1704), .Y(n2026) );
  CLKBUFX3 U1386 ( .A(n2023), .Y(n1700) );
  NAND2XL U1387 ( .A(n1626), .B(n1702), .Y(n2023) );
  CLKBUFX3 U1388 ( .A(n2018), .Y(n1697) );
  NAND2XL U1389 ( .A(n1626), .B(n1699), .Y(n2018) );
  CLKBUFX3 U1390 ( .A(n2157), .Y(n1715) );
  NAND2XL U1391 ( .A(n1614), .B(n1717), .Y(n2157) );
  CLKBUFX3 U1392 ( .A(n2190), .Y(n1723) );
  NAND2X1 U1393 ( .A(n1587), .B(n1724), .Y(n2190) );
  CLKBUFX3 U1394 ( .A(n2187), .Y(n1720) );
  NAND2XL U1395 ( .A(n1587), .B(n1721), .Y(n2187) );
  CLKBUFX3 U1396 ( .A(n2211), .Y(n1739) );
  CLKBUFX3 U1397 ( .A(n1480), .Y(n1737) );
  CLKBUFX3 U1398 ( .A(n2194), .Y(n1725) );
  NAND2XL U1399 ( .A(n1587), .B(n1726), .Y(n2194) );
  CLKBUFX3 U1400 ( .A(n2161), .Y(n1718) );
  NAND2XL U1401 ( .A(n1614), .B(n1719), .Y(n2161) );
  CLKBUFX3 U1402 ( .A(n1853), .Y(n1733) );
  CLKBUFX3 U1403 ( .A(n1808), .Y(n1689) );
  NAND3X1 U1404 ( .A(n1914), .B(n1915), .C(n1916), .Y(n1808) );
  CLKBUFX3 U1405 ( .A(n2619), .Y(n1767) );
  AND2X2 U1406 ( .A(n1918), .B(n1934), .Y(n1897) );
  AND2X2 U1407 ( .A(n1912), .B(n1954), .Y(n1890) );
  CLKBUFX3 U1408 ( .A(n1827), .Y(n1729) );
  NAND2X1 U1409 ( .A(state[1]), .B(n2503), .Y(n1827) );
  CLKBUFX3 U1410 ( .A(n1813), .Y(n1728) );
  NAND2X1 U1411 ( .A(n1994), .B(state[1]), .Y(n1813) );
  NAND3X2 U1412 ( .A(n1724), .B(n1847), .C(n2586), .Y(n2189) );
  NAND3X2 U1413 ( .A(n2081), .B(n1695), .C(n2618), .Y(n2007) );
  NAND3X2 U1414 ( .A(n1713), .B(n2394), .C(n2599), .Y(n2150) );
  NAND3X2 U1415 ( .A(n2599), .B(n1713), .C(n2395), .Y(n2146) );
  CLKBUFX3 U1416 ( .A(n2022), .Y(n1701) );
  NAND3X1 U1417 ( .A(n1841), .B(n1702), .C(n2618), .Y(n2022) );
  CLKBUFX3 U1418 ( .A(n2156), .Y(n1716) );
  NAND3X1 U1419 ( .A(n1842), .B(n1717), .C(n2599), .Y(n2156) );
  NAND2X2 U1420 ( .A(n2618), .B(n1704), .Y(n2028) );
  NAND2X2 U1421 ( .A(n2586), .B(n1721), .Y(n2188) );
  NAND2X2 U1422 ( .A(n2618), .B(n1706), .Y(n2015) );
  AND3X4 U1423 ( .A(n1695), .B(n2618), .C(n2080), .Y(n2010) );
  AND3X4 U1424 ( .A(n1702), .B(n1814), .C(n2618), .Y(n2025) );
  AND3X4 U1425 ( .A(n1717), .B(n2102), .C(n2599), .Y(n2159) );
  INVX3 U1426 ( .A(sort_stage[0]), .Y(n1830) );
  CLKBUFX3 U1427 ( .A(n2012), .Y(n1706) );
  OAI31XL U1428 ( .A0(n1838), .A1(n2132), .A2(n1822), .B0(n2084), .Y(n2012) );
  CLKBUFX3 U1429 ( .A(n2196), .Y(n1726) );
  OAI31XL U1430 ( .A0(n1847), .A1(n2459), .A2(n1729), .B0(n2257), .Y(n2196) );
  CLKBUFX3 U1431 ( .A(n2029), .Y(n1704) );
  OAI31XL U1432 ( .A0(n1814), .A1(n2117), .A2(n1822), .B0(n2084), .Y(n2029) );
  CLKBUFX3 U1433 ( .A(n2151), .Y(n1714) );
  OAI31XL U1434 ( .A0(n1838), .A1(n2396), .A2(n1728), .B0(n2258), .Y(n2151) );
  CLKBUFX3 U1435 ( .A(n2192), .Y(n1722) );
  NAND3XL U1436 ( .A(n1843), .B(n1724), .C(n2586), .Y(n2192) );
  CLKBUFX3 U1437 ( .A(n2017), .Y(n1698) );
  NAND3X1 U1438 ( .A(n2618), .B(n1699), .C(n2083), .Y(n2017) );
  CLKBUFX3 U1439 ( .A(n1826), .Y(n1730) );
  NAND2X1 U1440 ( .A(n2504), .B(state[0]), .Y(n1826) );
  CLKINVX1 U1441 ( .A(n1686), .Y(n2211) );
  NAND2X2 U1442 ( .A(n2586), .B(n1726), .Y(n2195) );
  NAND2X2 U1443 ( .A(n2599), .B(n1719), .Y(n2162) );
  NAND2X2 U1444 ( .A(n2599), .B(n1714), .Y(n2154) );
  CLKBUFX3 U1445 ( .A(n2163), .Y(n1719) );
  OAI31XL U1446 ( .A0(n2102), .A1(n2426), .A2(n1728), .B0(n2258), .Y(n2163) );
  NAND2BX1 U1447 ( .AN(gray_valid), .B(n1688), .Y(n1687) );
  CLKINVX1 U1448 ( .A(n1687), .Y(n1853) );
  CLKBUFX3 U1449 ( .A(n1807), .Y(n1693) );
  NAND3X1 U1450 ( .A(n1916), .B(n1914), .C(gray_data[1]), .Y(n1807) );
  CLKBUFX3 U1451 ( .A(n1812), .Y(n1694) );
  NAND3X1 U1452 ( .A(n1932), .B(n1915), .C(gray_data[0]), .Y(n1812) );
  CLKBUFX3 U1453 ( .A(n1810), .Y(n1692) );
  NAND3XL U1454 ( .A(n1916), .B(n1915), .C(gray_data[0]), .Y(n1810) );
  CLKBUFX3 U1455 ( .A(n1811), .Y(n1690) );
  NAND3X1 U1456 ( .A(n1932), .B(gray_data[1]), .C(gray_data[0]), .Y(n1811) );
  CLKBUFX3 U1457 ( .A(n1809), .Y(n1691) );
  NAND3XL U1458 ( .A(gray_data[1]), .B(n1914), .C(n1932), .Y(n1809) );
  NAND2BX1 U1459 ( .AN(\C4[0][4] ), .B(\C4[1][4] ), .Y(n1769) );
  OAI222XL U1460 ( .A0(\C4[0][5] ), .A1(n877), .B0(\C4[0][5] ), .B1(n1769), 
        .C0(n877), .C1(n1769), .Y(n1770) );
  OAI222XL U1461 ( .A0(\C4[1][6] ), .A1(n1770), .B0(n876), .B1(n1770), .C0(
        \C4[1][6] ), .C1(n876), .Y(n1781) );
  NAND2BX1 U1462 ( .AN(\C4[0][2] ), .B(\C4[1][2] ), .Y(n1773) );
  OAI22XL U1463 ( .A0(\C4[0][3] ), .A1(n881), .B0(\C4[0][3] ), .B1(n1773), .Y(
        n1779) );
  NOR2BX1 U1464 ( .AN(\C4[0][2] ), .B(\C4[1][2] ), .Y(n1771) );
  OA22X1 U1465 ( .A0(n1771), .A1(\C4[0][3] ), .B0(n1771), .B1(n881), .Y(n1775)
         );
  AOI21X1 U1466 ( .A0(\C4[0][1] ), .A1(n885), .B0(\C4[0][0] ), .Y(n1772) );
  AOI2BB2X1 U1467 ( .B0(n1772), .B1(\C4[1][0] ), .A0N(\C4[0][1] ), .A1N(n885), 
        .Y(n1774) );
  OAI22XL U1468 ( .A0(n1775), .A1(n1774), .B0(n1773), .B1(n881), .Y(n1778) );
  NOR2BX1 U1469 ( .AN(\C4[0][4] ), .B(\C4[1][4] ), .Y(n1776) );
  OAI22XL U1470 ( .A0(n1776), .A1(n877), .B0(\C4[0][5] ), .B1(n1776), .Y(n1777) );
  OAI221XL U1471 ( .A0(\C4[1][6] ), .A1(n876), .B0(n1779), .B1(n1778), .C0(
        n1777), .Y(n1780) );
  AO22X1 U1472 ( .A0(n889), .A1(\C4[0][7] ), .B0(n1781), .B1(n1780), .Y(n1782)
         );
  OAI21XL U1473 ( .A0(\C4[0][7] ), .A1(n889), .B0(n1782), .Y(N2784) );
  CLKINVX1 U1474 ( .A(reset), .Y(n2619) );
  NAND2X1 U1475 ( .A(n1783), .B(n1784), .Y(n2620) );
  MXI2X1 U1476 ( .A(n2557), .B(n1785), .S0(n1727), .Y(n1783) );
  NAND2X1 U1477 ( .A(n1787), .B(n1788), .Y(n2621) );
  MXI2X1 U1478 ( .A(n2548), .B(n1789), .S0(n1712), .Y(n1787) );
  NAND2X1 U1479 ( .A(n1791), .B(n1792), .Y(n2622) );
  MXI2X1 U1480 ( .A(n2539), .B(n1793), .S0(n1711), .Y(n1791) );
  NAND2X1 U1481 ( .A(n1795), .B(n1796), .Y(n2623) );
  MXI2X1 U1482 ( .A(n2530), .B(n1797), .S0(n1710), .Y(n1795) );
  NAND2X1 U1483 ( .A(n1799), .B(n1800), .Y(n2624) );
  MXI2X1 U1484 ( .A(n2521), .B(n1801), .S0(n1709), .Y(n1799) );
  NAND2X1 U1485 ( .A(n1803), .B(n1804), .Y(n2625) );
  MXI2X1 U1486 ( .A(n2511), .B(n1805), .S0(n1707), .Y(n1803) );
  CLKMX2X2 U1487 ( .A(N967), .B(CNT6[0]), .S0(n1693), .Y(n1477) );
  CLKMX2X2 U1488 ( .A(N968), .B(CNT6[1]), .S0(n1693), .Y(n1476) );
  CLKMX2X2 U1489 ( .A(N969), .B(CNT6[2]), .S0(n1693), .Y(n1475) );
  CLKMX2X2 U1490 ( .A(N970), .B(CNT6[3]), .S0(n1693), .Y(n1474) );
  CLKMX2X2 U1491 ( .A(N971), .B(CNT6[4]), .S0(n1693), .Y(n1473) );
  CLKMX2X2 U1492 ( .A(N972), .B(CNT6[5]), .S0(n1693), .Y(n1472) );
  CLKMX2X2 U1493 ( .A(N973), .B(CNT6[6]), .S0(n1693), .Y(n1471) );
  CLKMX2X2 U1494 ( .A(N974), .B(CNT6[7]), .S0(n1693), .Y(n1470) );
  CLKMX2X2 U1495 ( .A(N935), .B(CNT4[0]), .S0(n1689), .Y(n1469) );
  CLKMX2X2 U1496 ( .A(N936), .B(CNT4[1]), .S0(n1689), .Y(n1468) );
  CLKMX2X2 U1497 ( .A(N937), .B(CNT4[2]), .S0(n1689), .Y(n1467) );
  CLKMX2X2 U1498 ( .A(N938), .B(CNT4[3]), .S0(n1689), .Y(n1466) );
  CLKMX2X2 U1499 ( .A(N939), .B(CNT4[4]), .S0(n1689), .Y(n1465) );
  CLKMX2X2 U1500 ( .A(N940), .B(CNT4[5]), .S0(n1689), .Y(n1464) );
  CLKMX2X2 U1501 ( .A(N941), .B(CNT4[6]), .S0(n1689), .Y(n1463) );
  CLKMX2X2 U1502 ( .A(N942), .B(CNT4[7]), .S0(n1689), .Y(n1462) );
  CLKMX2X2 U1503 ( .A(N903), .B(CNT2[0]), .S0(n1691), .Y(n1461) );
  CLKMX2X2 U1504 ( .A(N904), .B(CNT2[1]), .S0(n1691), .Y(n1460) );
  CLKMX2X2 U1505 ( .A(N905), .B(CNT2[2]), .S0(n1691), .Y(n1459) );
  CLKMX2X2 U1506 ( .A(N906), .B(CNT2[3]), .S0(n1691), .Y(n1458) );
  CLKMX2X2 U1507 ( .A(N907), .B(CNT2[4]), .S0(n1691), .Y(n1457) );
  CLKMX2X2 U1508 ( .A(N908), .B(CNT2[5]), .S0(n1691), .Y(n1456) );
  CLKMX2X2 U1509 ( .A(N909), .B(CNT2[6]), .S0(n1691), .Y(n1455) );
  CLKMX2X2 U1510 ( .A(N910), .B(CNT2[7]), .S0(n1691), .Y(n1454) );
  CLKMX2X2 U1511 ( .A(N951), .B(CNT5[0]), .S0(n1692), .Y(n1453) );
  CLKMX2X2 U1512 ( .A(N952), .B(CNT5[1]), .S0(n1692), .Y(n1452) );
  CLKMX2X2 U1513 ( .A(N953), .B(CNT5[2]), .S0(n1692), .Y(n1451) );
  CLKMX2X2 U1514 ( .A(N954), .B(CNT5[3]), .S0(n1692), .Y(n1450) );
  CLKMX2X2 U1515 ( .A(N955), .B(CNT5[4]), .S0(n1692), .Y(n1449) );
  CLKMX2X2 U1516 ( .A(N956), .B(CNT5[5]), .S0(n1692), .Y(n1448) );
  CLKMX2X2 U1517 ( .A(N957), .B(CNT5[6]), .S0(n1692), .Y(n1447) );
  CLKMX2X2 U1518 ( .A(N958), .B(CNT5[7]), .S0(n1692), .Y(n1446) );
  CLKMX2X2 U1519 ( .A(N919), .B(CNT3[0]), .S0(n1690), .Y(n1445) );
  CLKMX2X2 U1520 ( .A(N920), .B(CNT3[1]), .S0(n1690), .Y(n1444) );
  CLKMX2X2 U1521 ( .A(N921), .B(CNT3[2]), .S0(n1690), .Y(n1443) );
  CLKMX2X2 U1522 ( .A(N922), .B(CNT3[3]), .S0(n1690), .Y(n1442) );
  CLKMX2X2 U1523 ( .A(N923), .B(CNT3[4]), .S0(n1690), .Y(n1441) );
  CLKMX2X2 U1524 ( .A(N924), .B(CNT3[5]), .S0(n1690), .Y(n1440) );
  CLKMX2X2 U1525 ( .A(N925), .B(CNT3[6]), .S0(n1690), .Y(n1439) );
  CLKMX2X2 U1526 ( .A(N926), .B(CNT3[7]), .S0(n1690), .Y(n1438) );
  CLKMX2X2 U1527 ( .A(N887), .B(CNT1[0]), .S0(n1694), .Y(n1437) );
  CLKMX2X2 U1528 ( .A(N888), .B(CNT1[1]), .S0(n1694), .Y(n1436) );
  CLKMX2X2 U1529 ( .A(N889), .B(CNT1[2]), .S0(n1694), .Y(n1435) );
  CLKMX2X2 U1530 ( .A(N890), .B(CNT1[3]), .S0(n1694), .Y(n1434) );
  CLKMX2X2 U1531 ( .A(N891), .B(CNT1[4]), .S0(n1694), .Y(n1433) );
  CLKMX2X2 U1532 ( .A(N892), .B(CNT1[5]), .S0(n1694), .Y(n1432) );
  CLKMX2X2 U1533 ( .A(N893), .B(CNT1[6]), .S0(n1694), .Y(n1431) );
  CLKMX2X2 U1534 ( .A(N894), .B(CNT1[7]), .S0(n1694), .Y(n1430) );
  OAI21XL U1535 ( .A0(n1814), .A1(n1815), .B0(n1816), .Y(n1428) );
  OAI21XL U1536 ( .A0(n1581), .A1(n1817), .B0(sort_stage[2]), .Y(n1816) );
  NAND2X1 U1537 ( .A(n1818), .B(n1819), .Y(n1427) );
  CLKMX2X2 U1538 ( .A(n1820), .B(n1580), .S0(n1821), .Y(n1818) );
  MXI2X1 U1539 ( .A(n1823), .B(n1583), .S0(n1821), .Y(n1425) );
  NOR2X1 U1540 ( .A(n1824), .B(n1825), .Y(n1823) );
  NAND2X1 U1541 ( .A(n1019), .B(n1730), .Y(n1424) );
  OAI21XL U1542 ( .A0(n1821), .A1(n1729), .B0(n1586), .Y(n1423) );
  NAND2X1 U1543 ( .A(n1587), .B(n1729), .Y(n1421) );
  MXI2X1 U1544 ( .A(n1829), .B(n1815), .S0(n1830), .Y(n1420) );
  MXI2X1 U1545 ( .A(n1831), .B(n1832), .S0(n1581), .Y(n1419) );
  OR2X1 U1546 ( .A(n1815), .B(n1830), .Y(n1832) );
  NAND2BX1 U1547 ( .AN(n1833), .B(n1829), .Y(n1815) );
  CLKINVX1 U1548 ( .A(n1817), .Y(n1831) );
  OAI21XL U1549 ( .A0(sort_stage[0]), .A1(n1833), .B0(n1829), .Y(n1817) );
  OR4X1 U1550 ( .A(n1834), .B(n1835), .C(n1836), .D(n1837), .Y(n1829) );
  OAI31XL U1551 ( .A0(n1838), .A1(n1729), .A2(n1587), .B0(n1821), .Y(n1837) );
  AND2X1 U1552 ( .A(n1839), .B(n1840), .Y(n1821) );
  AOI33X1 U1553 ( .A0(n1841), .A1(n1825), .A2(n2618), .B0(n1842), .B1(n1824), 
        .B2(n2599), .Y(n1840) );
  OAI21XL U1554 ( .A0(n1848), .A1(n1849), .B0(n1586), .Y(n1833) );
  MXI2X1 U1555 ( .A(n1850), .B(n1842), .S0(n1580), .Y(n1849) );
  NAND2X1 U1556 ( .A(state[1]), .B(n1847), .Y(n1850) );
  NOR2X1 U1557 ( .A(state[1]), .B(n1841), .Y(n1848) );
  OAI21XL U1558 ( .A0(n1017), .A1(n1825), .B0(n1819), .Y(n1418) );
  NAND4X1 U1559 ( .A(n1834), .B(sort_stage[0]), .C(sort_stage[1]), .D(
        sort_stage[2]), .Y(n1819) );
  AOI222XL U1560 ( .A0(N966), .A1(gray_valid), .B0(n1478), .B1(
        \symbol_value[3][7] ), .C0(n1734), .C1(\symbol_value[5][7] ), .Y(n1851) );
  CLKINVX1 U1561 ( .A(n1854), .Y(n1416) );
  AOI222XL U1562 ( .A0(n1855), .A1(\symbol_value[5][7] ), .B0(n1856), .B1(
        \symbol_value[4][7] ), .C0(N982), .C1(n1857), .Y(n1854) );
  CLKINVX1 U1563 ( .A(n1858), .Y(n1415) );
  AOI222XL U1564 ( .A0(\symbol_value[5][6] ), .A1(n1855), .B0(n1856), .B1(
        \symbol_value[4][6] ), .C0(N981), .C1(n1857), .Y(n1858) );
  AOI222XL U1565 ( .A0(N965), .A1(gray_valid), .B0(n1478), .B1(
        \symbol_value[3][6] ), .C0(\symbol_value[5][6] ), .C1(n1733), .Y(n1859) );
  AOI222XL U1566 ( .A0(N949), .A1(gray_valid), .B0(n1478), .B1(
        \symbol_value[4][6] ), .C0(\symbol_value[2][6] ), .C1(n1733), .Y(n1860) );
  AOI222XL U1567 ( .A0(N933), .A1(gray_valid), .B0(\symbol_value[1][6] ), .B1(
        n1732), .C0(n1734), .C1(\symbol_value[3][6] ), .Y(n1862) );
  AOI222XL U1568 ( .A0(N917), .A1(gray_valid), .B0(\symbol_value[2][6] ), .B1(
        n1478), .C0(\symbol_value[0][6] ), .C1(n1733), .Y(n1864) );
  CLKINVX1 U1569 ( .A(n1866), .Y(n1410) );
  AOI222XL U1570 ( .A0(n1867), .A1(\symbol_value[0][6] ), .B0(n1868), .B1(
        \symbol_value[1][6] ), .C0(N901), .C1(n1869), .Y(n1866) );
  AOI222XL U1571 ( .A0(N918), .A1(gray_valid), .B0(\symbol_value[2][7] ), .B1(
        n1731), .C0(\symbol_value[0][7] ), .C1(n1733), .Y(n1870) );
  CLKINVX1 U1572 ( .A(n1871), .Y(n1408) );
  AOI222XL U1573 ( .A0(n1867), .A1(\symbol_value[0][7] ), .B0(n1868), .B1(
        \symbol_value[1][7] ), .C0(N902), .C1(n1869), .Y(n1871) );
  CLKINVX1 U1574 ( .A(n1872), .Y(n1407) );
  AOI222XL U1575 ( .A0(n1867), .A1(\symbol_value[0][5] ), .B0(n1868), .B1(
        \symbol_value[1][5] ), .C0(N900), .C1(n1869), .Y(n1872) );
  AOI222XL U1576 ( .A0(N916), .A1(gray_valid), .B0(\symbol_value[2][5] ), .B1(
        n1732), .C0(\symbol_value[0][5] ), .C1(n1733), .Y(n1873) );
  AOI222XL U1577 ( .A0(N932), .A1(gray_valid), .B0(\symbol_value[1][5] ), .B1(
        n1732), .C0(n1734), .C1(\symbol_value[3][5] ), .Y(n1874) );
  AOI222XL U1578 ( .A0(N948), .A1(gray_valid), .B0(n1732), .B1(
        \symbol_value[4][5] ), .C0(\symbol_value[2][5] ), .C1(n1734), .Y(n1875) );
  AOI222XL U1579 ( .A0(N964), .A1(gray_valid), .B0(n1732), .B1(
        \symbol_value[3][5] ), .C0(n1734), .C1(\symbol_value[5][5] ), .Y(n1876) );
  CLKINVX1 U1580 ( .A(n1877), .Y(n1402) );
  AOI222XL U1581 ( .A0(n1855), .A1(\symbol_value[5][5] ), .B0(n1856), .B1(
        \symbol_value[4][5] ), .C0(N980), .C1(n1857), .Y(n1877) );
  CLKINVX1 U1582 ( .A(n1878), .Y(n1401) );
  AOI222XL U1583 ( .A0(n1855), .A1(\symbol_value[5][4] ), .B0(n1856), .B1(
        \symbol_value[4][4] ), .C0(N979), .C1(n1857), .Y(n1878) );
  AOI222XL U1584 ( .A0(N963), .A1(gray_valid), .B0(n1732), .B1(
        \symbol_value[3][4] ), .C0(n1734), .C1(\symbol_value[5][4] ), .Y(n1879) );
  AOI222XL U1585 ( .A0(N947), .A1(gray_valid), .B0(n1732), .B1(
        \symbol_value[4][4] ), .C0(\symbol_value[2][4] ), .C1(n1734), .Y(n1880) );
  AOI222XL U1586 ( .A0(N931), .A1(gray_valid), .B0(\symbol_value[1][4] ), .B1(
        n1732), .C0(n1734), .C1(\symbol_value[3][4] ), .Y(n1881) );
  AOI222XL U1587 ( .A0(N915), .A1(gray_valid), .B0(\symbol_value[2][4] ), .B1(
        n1732), .C0(\symbol_value[0][4] ), .C1(n1734), .Y(n1882) );
  AOI222XL U1588 ( .A0(N934), .A1(gray_valid), .B0(\symbol_value[1][7] ), .B1(
        n1732), .C0(n1734), .C1(\symbol_value[3][7] ), .Y(n1883) );
  AOI222XL U1589 ( .A0(N950), .A1(gray_valid), .B0(n1732), .B1(
        \symbol_value[4][7] ), .C0(\symbol_value[2][7] ), .C1(n1734), .Y(n1884) );
  OAI222XL U1590 ( .A0(n1885), .A1(n1493), .B0(n1886), .B1(n1482), .C0(n1887), 
        .C1(n1553), .Y(n1394) );
  OAI222XL U1591 ( .A0(n1553), .A1(n1888), .B0(n1889), .B1(n1655), .C0(n1890), 
        .C1(n1493), .Y(n1393) );
  OAI222XL U1592 ( .A0(n1892), .A1(n1520), .B0(n1553), .B1(n1893), .C0(n1894), 
        .C1(n1482), .Y(n1391) );
  OAI222XL U1593 ( .A0(n1482), .A1(n1895), .B0(n1896), .B1(n1651), .C0(n1897), 
        .C1(n1520), .Y(n1390) );
  OAI222XL U1594 ( .A0(n1885), .A1(n1494), .B0(n1886), .B1(n1486), .C0(n1887), 
        .C1(n1554), .Y(n1388) );
  OAI222XL U1595 ( .A0(n1888), .A1(n1554), .B0(n1889), .B1(n1656), .C0(n1890), 
        .C1(n1494), .Y(n1387) );
  OAI222XL U1596 ( .A0(n1892), .A1(n1519), .B0(n1893), .B1(n1554), .C0(n1894), 
        .C1(n1486), .Y(n1385) );
  OAI222XL U1597 ( .A0(n1895), .A1(n1486), .B0(n1896), .B1(n1650), .C0(n1897), 
        .C1(n1519), .Y(n1384) );
  OAI222XL U1598 ( .A0(n1885), .A1(n1495), .B0(n1886), .B1(n1485), .C0(n1887), 
        .C1(n1555), .Y(n1382) );
  OAI222XL U1599 ( .A0(n1888), .A1(n1555), .B0(n1889), .B1(n1657), .C0(n1890), 
        .C1(n1495), .Y(n1381) );
  OAI222XL U1600 ( .A0(n1892), .A1(n1518), .B0(n1893), .B1(n1555), .C0(n1894), 
        .C1(n1485), .Y(n1379) );
  OAI222XL U1601 ( .A0(n1895), .A1(n1485), .B0(n1896), .B1(n1649), .C0(n1897), 
        .C1(n1518), .Y(n1378) );
  OAI222XL U1602 ( .A0(n1885), .A1(n1521), .B0(n1886), .B1(n1484), .C0(n1887), 
        .C1(n1557), .Y(n1376) );
  OAI222XL U1603 ( .A0(n1888), .A1(n1557), .B0(n1889), .B1(n1658), .C0(n1890), 
        .C1(n1521), .Y(n1375) );
  OAI222XL U1604 ( .A0(n1892), .A1(n1517), .B0(n1893), .B1(n1557), .C0(n1894), 
        .C1(n1484), .Y(n1373) );
  OAI222XL U1605 ( .A0(n1895), .A1(n1484), .B0(n1896), .B1(n1648), .C0(n1897), 
        .C1(n1517), .Y(n1372) );
  OAI222XL U1606 ( .A0(n1885), .A1(n1496), .B0(n1886), .B1(n1483), .C0(n1887), 
        .C1(n1556), .Y(n1370) );
  OAI222XL U1607 ( .A0(n1888), .A1(n1556), .B0(n1889), .B1(n1659), .C0(n1890), 
        .C1(n1496), .Y(n1369) );
  OAI222XL U1608 ( .A0(n1892), .A1(n1516), .B0(n1893), .B1(n1556), .C0(n1894), 
        .C1(n1483), .Y(n1367) );
  OAI222XL U1609 ( .A0(n1895), .A1(n1483), .B0(n1896), .B1(n1647), .C0(n1897), 
        .C1(n1516), .Y(n1366) );
  OAI222XL U1610 ( .A0(n1885), .A1(n1564), .B0(n1886), .B1(n1479), .C0(n1887), 
        .C1(n1522), .Y(n1364) );
  NAND2X1 U1611 ( .A(n1887), .B(n1830), .Y(n1886) );
  NAND2X1 U1612 ( .A(n1887), .B(sort_stage[0]), .Y(n1885) );
  OAI222XL U1613 ( .A0(n1888), .A1(n1522), .B0(n1889), .B1(n1684), .C0(n1890), 
        .C1(n1564), .Y(n1363) );
  NAND2X1 U1614 ( .A(n1890), .B(n1830), .Y(n1889) );
  NAND2X1 U1615 ( .A(n1890), .B(sort_stage[0]), .Y(n1888) );
  OAI222XL U1616 ( .A0(n1892), .A1(n1487), .B0(n1893), .B1(n1522), .C0(n1894), 
        .C1(n1479), .Y(n1361) );
  NAND2X1 U1617 ( .A(n1894), .B(n1830), .Y(n1893) );
  NAND2X1 U1618 ( .A(n1894), .B(sort_stage[0]), .Y(n1892) );
  OAI222XL U1619 ( .A0(n1895), .A1(n1479), .B0(n1896), .B1(n1646), .C0(n1897), 
        .C1(n1487), .Y(n1360) );
  NAND2X1 U1620 ( .A(n1897), .B(n1830), .Y(n1896) );
  NAND2X1 U1621 ( .A(n1897), .B(sort_stage[0]), .Y(n1895) );
  AOI222XL U1622 ( .A0(N946), .A1(gray_valid), .B0(n1732), .B1(
        \symbol_value[4][3] ), .C0(\symbol_value[2][3] ), .C1(n1734), .Y(n1899) );
  AOI222XL U1623 ( .A0(N962), .A1(gray_valid), .B0(n1732), .B1(
        \symbol_value[3][3] ), .C0(n1733), .C1(\symbol_value[5][3] ), .Y(n1900) );
  AOI222XL U1624 ( .A0(N961), .A1(gray_valid), .B0(n1732), .B1(
        \symbol_value[3][2] ), .C0(n1853), .C1(\symbol_value[5][2] ), .Y(n1901) );
  AOI222XL U1625 ( .A0(N945), .A1(gray_valid), .B0(n1731), .B1(
        \symbol_value[4][2] ), .C0(\symbol_value[2][2] ), .C1(n1733), .Y(n1902) );
  AOI222XL U1626 ( .A0(N929), .A1(gray_valid), .B0(\symbol_value[1][2] ), .B1(
        n1731), .C0(n1734), .C1(\symbol_value[3][2] ), .Y(n1903) );
  AOI222XL U1627 ( .A0(N913), .A1(gray_valid), .B0(\symbol_value[2][2] ), .B1(
        n1731), .C0(\symbol_value[0][2] ), .C1(n1733), .Y(n1904) );
  AOI222XL U1628 ( .A0(N914), .A1(gray_valid), .B0(\symbol_value[2][3] ), .B1(
        n1731), .C0(\symbol_value[0][3] ), .C1(n1733), .Y(n1905) );
  AOI222XL U1629 ( .A0(N930), .A1(gray_valid), .B0(\symbol_value[1][3] ), .B1(
        n1731), .C0(n1733), .C1(\symbol_value[3][3] ), .Y(n1906) );
  AOI222XL U1630 ( .A0(N928), .A1(gray_valid), .B0(\symbol_value[1][1] ), .B1(
        n1731), .C0(n1734), .C1(\symbol_value[3][1] ), .Y(n1907) );
  AOI222XL U1631 ( .A0(N912), .A1(gray_valid), .B0(\symbol_value[2][1] ), .B1(
        n1731), .C0(\symbol_value[0][1] ), .C1(n1733), .Y(n1908) );
  CLKINVX1 U1632 ( .A(n1909), .Y(n1348) );
  AOI222XL U1633 ( .A0(n1867), .A1(\symbol_value[0][1] ), .B0(n1868), .B1(
        \symbol_value[1][1] ), .C0(N896), .C1(n1869), .Y(n1909) );
  AOI222XL U1634 ( .A0(N944), .A1(gray_valid), .B0(n1731), .B1(
        \symbol_value[4][1] ), .C0(\symbol_value[2][1] ), .C1(n1733), .Y(n1910) );
  MXI2X1 U1635 ( .A(n1911), .B(n1618), .S0(n1861), .Y(n1346) );
  AOI222XL U1636 ( .A0(N943), .A1(gray_valid), .B0(n1731), .B1(
        \symbol_value[4][0] ), .C0(\symbol_value[2][0] ), .C1(n1733), .Y(n1911) );
  MXI2X1 U1637 ( .A(n1917), .B(n1606), .S0(n1863), .Y(n1345) );
  OAI221XL U1638 ( .A0(n1919), .A1(n1920), .B0(\symbol_value[2][7] ), .B1(
        n1625), .C0(n1830), .Y(n1913) );
  NOR2X1 U1639 ( .A(\symbol_value[3][7] ), .B(n1621), .Y(n1920) );
  AOI32X1 U1640 ( .A0(n1921), .A1(n1922), .A2(n1923), .B0(n1924), .B1(n1925), 
        .Y(n1919) );
  OAI21XL U1641 ( .A0(n1926), .A1(\symbol_value[2][6] ), .B0(n1624), .Y(n1925)
         );
  NAND2X1 U1642 ( .A(n1926), .B(\symbol_value[2][6] ), .Y(n1924) );
  AOI32X1 U1643 ( .A0(\symbol_value[3][4] ), .A1(n1541), .A2(n1922), .B0(n1592), .B1(\symbol_value[3][5] ), .Y(n1926) );
  AOI2BB2X1 U1644 ( .B0(\symbol_value[2][6] ), .B1(n1624), .A0N(n1541), .A1N(
        \symbol_value[3][4] ), .Y(n1923) );
  NAND2X1 U1645 ( .A(\symbol_value[2][5] ), .B(n1543), .Y(n1922) );
  OAI211X1 U1646 ( .A0(n1540), .A1(n1927), .B0(n1928), .C0(n1929), .Y(n1921)
         );
  AO21X1 U1647 ( .A0(n1540), .A1(n1927), .B0(\symbol_value[2][3] ), .Y(n1929)
         );
  OAI222XL U1648 ( .A0(\symbol_value[3][3] ), .A1(n1538), .B0(
        \symbol_value[3][2] ), .B1(n1605), .C0(n1930), .C1(n1931), .Y(n1928)
         );
  NOR2X1 U1649 ( .A(\symbol_value[2][1] ), .B(n1544), .Y(n1931) );
  AOI211X1 U1650 ( .A0(\symbol_value[2][1] ), .A1(n1544), .B0(n1618), .C0(
        \symbol_value[2][0] ), .Y(n1930) );
  NAND2X1 U1651 ( .A(\symbol_value[3][2] ), .B(n1605), .Y(n1927) );
  AOI222XL U1652 ( .A0(N927), .A1(gray_valid), .B0(\symbol_value[1][0] ), .B1(
        n1731), .C0(\symbol_value[3][0] ), .C1(n1733), .Y(n1917) );
  MXI2X1 U1653 ( .A(n1933), .B(n1654), .S0(n1865), .Y(n1344) );
  OAI211X1 U1654 ( .A0(\symbol_value[0][7] ), .A1(n1620), .B0(n1935), .C0(
        n1830), .Y(n1934) );
  OA21XL U1655 ( .A0(n1830), .A1(n1936), .B0(n1834), .Y(n1918) );
  OAI22XL U1656 ( .A0(\symbol_value[1][7] ), .A1(n1621), .B0(n1937), .B1(n1938), .Y(n1936) );
  NOR2X1 U1657 ( .A(\symbol_value[2][7] ), .B(n1620), .Y(n1938) );
  AOI32X1 U1658 ( .A0(n1939), .A1(n1940), .A2(n1941), .B0(n1942), .B1(n1943), 
        .Y(n1937) );
  OAI21XL U1659 ( .A0(n1944), .A1(\symbol_value[1][6] ), .B0(n1622), .Y(n1943)
         );
  NAND2X1 U1660 ( .A(n1944), .B(\symbol_value[1][6] ), .Y(n1942) );
  AOI32X1 U1661 ( .A0(\symbol_value[2][4] ), .A1(n1539), .A2(n1940), .B0(n1604), .B1(\symbol_value[2][5] ), .Y(n1944) );
  AOI2BB2X1 U1662 ( .B0(\symbol_value[1][6] ), .B1(n1622), .A0N(n1539), .A1N(
        \symbol_value[2][4] ), .Y(n1941) );
  NAND2X1 U1663 ( .A(\symbol_value[1][5] ), .B(n1592), .Y(n1940) );
  OAI211X1 U1664 ( .A0(n1538), .A1(n1945), .B0(n1946), .C0(n1947), .Y(n1939)
         );
  AO21X1 U1665 ( .A0(n1538), .A1(n1945), .B0(\symbol_value[1][3] ), .Y(n1947)
         );
  OAI222XL U1666 ( .A0(\symbol_value[2][3] ), .A1(n1588), .B0(
        \symbol_value[2][2] ), .B1(n1527), .C0(n1948), .C1(n1949), .Y(n1946)
         );
  NOR2X1 U1667 ( .A(\symbol_value[1][1] ), .B(n1531), .Y(n1949) );
  AOI211X1 U1668 ( .A0(\symbol_value[1][1] ), .A1(n1531), .B0(n1606), .C0(
        \symbol_value[1][0] ), .Y(n1948) );
  NAND2X1 U1669 ( .A(\symbol_value[2][2] ), .B(n1527), .Y(n1945) );
  AOI222XL U1670 ( .A0(N911), .A1(gray_valid), .B0(\symbol_value[2][0] ), .B1(
        n1731), .C0(\symbol_value[0][0] ), .C1(n1733), .Y(n1933) );
  MXI2X1 U1671 ( .A(n1951), .B(n1608), .S0(n1852), .Y(n1342) );
  AOI222XL U1672 ( .A0(N959), .A1(gray_valid), .B0(\symbol_value[3][0] ), .B1(
        n1731), .C0(n1853), .C1(\symbol_value[5][0] ), .Y(n1951) );
  OAI211X1 U1673 ( .A0(\symbol_value[4][7] ), .A1(n1623), .B0(n1955), .C0(
        n1830), .Y(n1954) );
  OA21XL U1674 ( .A0(n1830), .A1(n1956), .B0(n1834), .Y(n1912) );
  OAI22XL U1675 ( .A0(\symbol_value[3][7] ), .A1(n1609), .B0(n1957), .B1(n1958), .Y(n1956) );
  NOR2X1 U1676 ( .A(\symbol_value[4][7] ), .B(n1625), .Y(n1958) );
  AOI32X1 U1677 ( .A0(n1959), .A1(n1960), .A2(n1961), .B0(n1962), .B1(n1963), 
        .Y(n1957) );
  OAI21XL U1678 ( .A0(n1964), .A1(\symbol_value[3][6] ), .B0(n1529), .Y(n1963)
         );
  NAND2X1 U1679 ( .A(n1964), .B(\symbol_value[3][6] ), .Y(n1962) );
  AOI32X1 U1680 ( .A0(\symbol_value[4][4] ), .A1(n1611), .A2(n1960), .B0(n1543), .B1(\symbol_value[4][5] ), .Y(n1964) );
  AOI2BB2X1 U1681 ( .B0(\symbol_value[3][6] ), .B1(n1529), .A0N(n1611), .A1N(
        \symbol_value[4][4] ), .Y(n1961) );
  NAND2X1 U1682 ( .A(\symbol_value[3][5] ), .B(n1530), .Y(n1960) );
  OAI211X1 U1683 ( .A0(n1965), .A1(n1591), .B0(n1966), .C0(n1967), .Y(n1959)
         );
  AO21X1 U1684 ( .A0(n1591), .A1(n1965), .B0(\symbol_value[3][3] ), .Y(n1967)
         );
  OAI222XL U1685 ( .A0(\symbol_value[4][3] ), .A1(n1540), .B0(
        \symbol_value[4][2] ), .B1(n1612), .C0(n1968), .C1(n1969), .Y(n1966)
         );
  NOR2X1 U1686 ( .A(\symbol_value[3][1] ), .B(n1528), .Y(n1969) );
  AOI211X1 U1687 ( .A0(\symbol_value[3][1] ), .A1(n1528), .B0(n1608), .C0(
        \symbol_value[3][0] ), .Y(n1968) );
  NAND2X1 U1688 ( .A(\symbol_value[4][2] ), .B(n1612), .Y(n1965) );
  AOI222XL U1689 ( .A0(N960), .A1(gray_valid), .B0(n1731), .B1(
        \symbol_value[3][1] ), .C0(n1734), .C1(\symbol_value[5][1] ), .Y(n1953) );
  CLKINVX1 U1690 ( .A(n1970), .Y(n1339) );
  AOI222XL U1691 ( .A0(n1855), .A1(\symbol_value[5][1] ), .B0(n1856), .B1(
        \symbol_value[4][1] ), .C0(N976), .C1(n1857), .Y(n1970) );
  CLKINVX1 U1692 ( .A(n1971), .Y(n1338) );
  AOI222XL U1693 ( .A0(n1867), .A1(\symbol_value[0][3] ), .B0(n1868), .B1(
        \symbol_value[1][3] ), .C0(N898), .C1(n1869), .Y(n1971) );
  CLKINVX1 U1694 ( .A(n1972), .Y(n1337) );
  AOI222XL U1695 ( .A0(n1867), .A1(\symbol_value[0][2] ), .B0(n1868), .B1(
        \symbol_value[1][2] ), .C0(N897), .C1(n1869), .Y(n1972) );
  CLKINVX1 U1696 ( .A(n1973), .Y(n1336) );
  AOI222XL U1697 ( .A0(n1855), .A1(\symbol_value[5][2] ), .B0(n1856), .B1(
        \symbol_value[4][2] ), .C0(N977), .C1(n1857), .Y(n1973) );
  CLKINVX1 U1698 ( .A(n1974), .Y(n1335) );
  AOI222XL U1699 ( .A0(n1855), .A1(\symbol_value[5][3] ), .B0(n1856), .B1(
        \symbol_value[4][3] ), .C0(N978), .C1(n1857), .Y(n1974) );
  NOR2X1 U1700 ( .A(\symbol_value[4][7] ), .B(n1623), .Y(n1976) );
  CLKINVX1 U1701 ( .A(n1955), .Y(n1975) );
  OAI21XL U1702 ( .A0(\symbol_value[5][7] ), .A1(n1609), .B0(n1977), .Y(n1955)
         );
  OAI32X1 U1703 ( .A0(n1978), .A1(n1979), .A2(n1980), .B0(n1981), .B1(n1982), 
        .Y(n1977) );
  AND2X1 U1704 ( .A(n1983), .B(\symbol_value[4][6] ), .Y(n1982) );
  AOI2BB1X1 U1705 ( .A0N(n1983), .A1N(\symbol_value[4][6] ), .B0(
        \symbol_value[5][6] ), .Y(n1981) );
  AOI32X1 U1706 ( .A0(\symbol_value[5][4] ), .A1(n1593), .A2(n1984), .B0(n1530), .B1(\symbol_value[5][5] ), .Y(n1983) );
  CLKINVX1 U1707 ( .A(n1979), .Y(n1984) );
  AOI211X1 U1708 ( .A0(\symbol_value[5][3] ), .A1(n1985), .B0(n1986), .C0(
        n1987), .Y(n1980) );
  AOI222XL U1709 ( .A0(n1988), .A1(n1989), .B0(\symbol_value[4][2] ), .B1(
        n1545), .C0(\symbol_value[4][3] ), .C1(n1619), .Y(n1987) );
  OAI211X1 U1710 ( .A0(\symbol_value[5][1] ), .A1(n1528), .B0(n1608), .C0(
        \symbol_value[5][0] ), .Y(n1989) );
  NAND2X1 U1711 ( .A(\symbol_value[5][1] ), .B(n1528), .Y(n1988) );
  OA21XL U1712 ( .A0(n1985), .A1(\symbol_value[5][3] ), .B0(n1591), .Y(n1986)
         );
  NOR2X1 U1713 ( .A(n1545), .B(\symbol_value[4][2] ), .Y(n1985) );
  NOR2X1 U1714 ( .A(n1530), .B(\symbol_value[5][5] ), .Y(n1979) );
  OAI22XL U1715 ( .A0(\symbol_value[5][6] ), .A1(n1529), .B0(
        \symbol_value[5][4] ), .B1(n1593), .Y(n1978) );
  CLKINVX1 U1716 ( .A(gray_data[0]), .Y(n1914) );
  NOR4BBX1 U1717 ( .AN(gray_data[2]), .BN(n1990), .C(gray_data[3]), .D(n1768), 
        .Y(n1916) );
  CLKINVX1 U1718 ( .A(n1991), .Y(n1334) );
  AOI222XL U1719 ( .A0(n1867), .A1(\symbol_value[0][4] ), .B0(n1868), .B1(
        \symbol_value[1][4] ), .C0(N899), .C1(n1869), .Y(n1991) );
  AND2X1 U1720 ( .A(n1994), .B(n1583), .Y(n1834) );
  NOR2X1 U1721 ( .A(\symbol_value[0][7] ), .B(n1620), .Y(n1993) );
  CLKINVX1 U1722 ( .A(n1935), .Y(n1992) );
  OAI21XL U1723 ( .A0(\symbol_value[1][7] ), .A1(n1610), .B0(n1995), .Y(n1935)
         );
  OAI32X1 U1724 ( .A0(n1996), .A1(n1997), .A2(n1998), .B0(n1999), .B1(n2000), 
        .Y(n1995) );
  NOR2X1 U1725 ( .A(n1542), .B(n2001), .Y(n2000) );
  AOI21X1 U1726 ( .A0(n1542), .A1(n2001), .B0(\symbol_value[1][6] ), .Y(n1999)
         );
  OAI32X1 U1727 ( .A0(n1539), .A1(\symbol_value[0][4] ), .A2(n1997), .B0(
        \symbol_value[0][5] ), .B1(n1604), .Y(n2001) );
  AOI221XL U1728 ( .A0(n1616), .A1(n2002), .B0(n2003), .B1(
        \symbol_value[1][3] ), .C0(n2004), .Y(n1998) );
  AOI222XL U1729 ( .A0(n2005), .A1(n2006), .B0(\symbol_value[0][2] ), .B1(
        n1527), .C0(\symbol_value[0][3] ), .C1(n1588), .Y(n2004) );
  OAI211X1 U1730 ( .A0(\symbol_value[1][1] ), .A1(n1535), .B0(n1596), .C0(
        \symbol_value[1][0] ), .Y(n2006) );
  NAND2X1 U1731 ( .A(\symbol_value[1][1] ), .B(n1535), .Y(n2005) );
  NAND2BX1 U1732 ( .AN(n2003), .B(n1588), .Y(n2002) );
  NOR2X1 U1733 ( .A(n1527), .B(\symbol_value[0][2] ), .Y(n2003) );
  NOR2X1 U1734 ( .A(n1597), .B(\symbol_value[1][5] ), .Y(n1997) );
  OAI22XL U1735 ( .A0(\symbol_value[1][6] ), .A1(n1542), .B0(
        \symbol_value[1][4] ), .B1(n1615), .Y(n1996) );
  CLKINVX1 U1736 ( .A(gray_data[1]), .Y(n1915) );
  NOR4BX1 U1737 ( .AN(n1990), .B(gray_data[2]), .C(gray_data[3]), .D(n1768), 
        .Y(n1932) );
  NOR4X1 U1738 ( .A(gray_data[7]), .B(gray_data[6]), .C(gray_data[5]), .D(
        gray_data[4]), .Y(n1990) );
  OAI221XL U1739 ( .A0(n1015), .A1(n2007), .B0(n1016), .B1(n1695), .C0(n2009), 
        .Y(n1333) );
  AOI22X1 U1740 ( .A0(n2010), .A1(n1579), .B0(n2011), .B1(\symbol_value[3][0] ), .Y(n2009) );
  OAI21XL U1741 ( .A0(n1015), .A1(n1706), .B0(n2013), .Y(n1332) );
  AOI2BB2X1 U1742 ( .B0(N1143), .B1(n1705), .A0N(n2015), .A1N(n1016), .Y(n2013) );
  OAI221XL U1743 ( .A0(n1012), .A1(n2007), .B0(n1013), .B1(n1695), .C0(n2016), 
        .Y(n1331) );
  AOI22X1 U1744 ( .A0(n2010), .A1(n1589), .B0(n2011), .B1(\symbol_value[3][7] ), .Y(n2016) );
  OAI221XL U1745 ( .A0(n1010), .A1(n1698), .B0(n1621), .B1(n1697), .C0(n2019), 
        .Y(n1330) );
  AOI2BB2X1 U1746 ( .B0(n1696), .B1(\C1[3][7] ), .A0N(n1699), .A1N(n1011), .Y(
        n2019) );
  OAI221XL U1747 ( .A0(n1009), .A1(n1701), .B0(n1620), .B1(n1700), .C0(n2024), 
        .Y(n1329) );
  AOI2BB2X1 U1748 ( .B0(n2025), .B1(n1589), .A0N(n1010), .A1N(n1702), .Y(n2024) );
  OAI222XL U1749 ( .A0(n1610), .A1(n1703), .B0(n1010), .B1(n2028), .C0(n1009), 
        .C1(n1704), .Y(n1328) );
  OAI221XL U1750 ( .A0(n1007), .A1(n1701), .B0(n1654), .B1(n1700), .C0(n2030), 
        .Y(n1327) );
  AOI2BB2X1 U1751 ( .B0(n2025), .B1(n1579), .A0N(n1008), .A1N(n1702), .Y(n2030) );
  OAI222XL U1752 ( .A0(n1596), .A1(n1703), .B0(n1008), .B1(n2028), .C0(n1007), 
        .C1(n1704), .Y(n1326) );
  OAI221XL U1753 ( .A0(n1008), .A1(n1698), .B0(n1606), .B1(n1697), .C0(n2031), 
        .Y(n1325) );
  AOI2BB2X1 U1754 ( .B0(n1696), .B1(\C1[3][0] ), .A0N(n1699), .A1N(n1014), .Y(
        n2031) );
  OAI221XL U1755 ( .A0(n1004), .A1(n1698), .B0(n1622), .B1(n1697), .C0(n2032), 
        .Y(n1324) );
  AOI2BB2X1 U1756 ( .B0(n1696), .B1(\C1[3][6] ), .A0N(n1699), .A1N(n1006), .Y(
        n2032) );
  OAI221XL U1757 ( .A0(n1003), .A1(n1701), .B0(n1652), .B1(n1700), .C0(n2033), 
        .Y(n1323) );
  AOI2BB2X1 U1758 ( .B0(n2025), .B1(n1590), .A0N(n1004), .A1N(n1702), .Y(n2033) );
  OAI222XL U1759 ( .A0(n1542), .A1(n1703), .B0(n1004), .B1(n2028), .C0(n1003), 
        .C1(n1704), .Y(n1322) );
  OAI221XL U1760 ( .A0(n1002), .A1(n2007), .B0(n1005), .B1(n1695), .C0(n2034), 
        .Y(n1321) );
  AOI22X1 U1761 ( .A0(n2010), .A1(n1590), .B0(n2011), .B1(\symbol_value[3][6] ), .Y(n2034) );
  OAI21XL U1762 ( .A0(n1002), .A1(n1706), .B0(n2035), .Y(n1320) );
  AOI2BB2X1 U1763 ( .B0(N1149), .B1(n1705), .A0N(n2015), .A1N(n1005), .Y(n2035) );
  OAI221XL U1764 ( .A0(n999), .A1(n1698), .B0(n1592), .B1(n1697), .C0(n2036), 
        .Y(n1319) );
  AOI2BB2X1 U1765 ( .B0(n1696), .B1(\C1[3][5] ), .A0N(n1699), .A1N(n1001), .Y(
        n2036) );
  OAI221XL U1766 ( .A0(n998), .A1(n1701), .B0(n1604), .B1(n1700), .C0(n2037), 
        .Y(n1318) );
  AOI2BB2X1 U1767 ( .B0(n2025), .B1(n1577), .A0N(n999), .A1N(n1702), .Y(n2037)
         );
  OAI222XL U1768 ( .A0(n1597), .A1(n1703), .B0(n999), .B1(n2028), .C0(n998), 
        .C1(n1704), .Y(n1317) );
  OAI221XL U1769 ( .A0(n997), .A1(n2007), .B0(n1000), .B1(n1695), .C0(n2038), 
        .Y(n1316) );
  AOI22X1 U1770 ( .A0(n2010), .A1(n1577), .B0(n2011), .B1(\symbol_value[3][5] ), .Y(n2038) );
  OAI21XL U1771 ( .A0(n997), .A1(n1706), .B0(n2039), .Y(n1315) );
  AOI2BB2X1 U1772 ( .B0(N1148), .B1(n1705), .A0N(n2015), .A1N(n1000), .Y(n2039) );
  OAI221XL U1773 ( .A0(n994), .A1(n1698), .B0(n1541), .B1(n1697), .C0(n2040), 
        .Y(n1314) );
  AOI2BB2X1 U1774 ( .B0(n1696), .B1(\C1[3][4] ), .A0N(n1699), .A1N(n996), .Y(
        n2040) );
  OAI221XL U1775 ( .A0(n993), .A1(n1701), .B0(n1539), .B1(n1700), .C0(n2041), 
        .Y(n1313) );
  AOI2BB2X1 U1776 ( .B0(n2025), .B1(n1525), .A0N(n994), .A1N(n1702), .Y(n2041)
         );
  OAI222XL U1777 ( .A0(n1615), .A1(n1703), .B0(n994), .B1(n2028), .C0(n993), 
        .C1(n1704), .Y(n1312) );
  OAI221XL U1778 ( .A0(n992), .A1(n2007), .B0(n995), .B1(n1695), .C0(n2042), 
        .Y(n1311) );
  AOI22X1 U1779 ( .A0(n2010), .A1(n1525), .B0(n2011), .B1(\symbol_value[3][4] ), .Y(n2042) );
  OAI21XL U1780 ( .A0(n992), .A1(n1706), .B0(n2043), .Y(n1310) );
  AOI2BB2X1 U1781 ( .B0(N1147), .B1(n1705), .A0N(n2015), .A1N(n995), .Y(n2043)
         );
  OAI221XL U1782 ( .A0(n989), .A1(n1698), .B0(n1538), .B1(n1697), .C0(n2044), 
        .Y(n1309) );
  AOI2BB2X1 U1783 ( .B0(n1696), .B1(\C1[3][3] ), .A0N(n1699), .A1N(n991), .Y(
        n2044) );
  OAI221XL U1784 ( .A0(n988), .A1(n1701), .B0(n1588), .B1(n1700), .C0(n2045), 
        .Y(n1308) );
  AOI2BB2X1 U1785 ( .B0(n2025), .B1(n1524), .A0N(n989), .A1N(n1702), .Y(n2045)
         );
  OAI222XL U1786 ( .A0(n1616), .A1(n1703), .B0(n989), .B1(n2028), .C0(n988), 
        .C1(n1704), .Y(n1307) );
  OAI221XL U1787 ( .A0(n987), .A1(n2007), .B0(n990), .B1(n1695), .C0(n2046), 
        .Y(n1306) );
  AOI22X1 U1788 ( .A0(n2010), .A1(n1524), .B0(n2011), .B1(\symbol_value[3][3] ), .Y(n2046) );
  OAI21XL U1789 ( .A0(n987), .A1(n1706), .B0(n2047), .Y(n1305) );
  AOI2BB2X1 U1790 ( .B0(N1146), .B1(n1705), .A0N(n2015), .A1N(n990), .Y(n2047)
         );
  OAI221XL U1791 ( .A0(n984), .A1(n1698), .B0(n1605), .B1(n1697), .C0(n2048), 
        .Y(n1304) );
  AOI2BB2X1 U1792 ( .B0(n1696), .B1(\C1[3][2] ), .A0N(n1699), .A1N(n986), .Y(
        n2048) );
  OAI221XL U1793 ( .A0(n983), .A1(n1701), .B0(n1527), .B1(n1700), .C0(n2049), 
        .Y(n1303) );
  AOI2BB2X1 U1794 ( .B0(n2025), .B1(n1578), .A0N(n984), .A1N(n1702), .Y(n2049)
         );
  OAI222XL U1795 ( .A0(n1639), .A1(n1703), .B0(n984), .B1(n2028), .C0(n983), 
        .C1(n1704), .Y(n1302) );
  OAI221XL U1796 ( .A0(n982), .A1(n2007), .B0(n985), .B1(n1695), .C0(n2050), 
        .Y(n1301) );
  AOI22X1 U1797 ( .A0(n2010), .A1(n1578), .B0(n2011), .B1(\symbol_value[3][2] ), .Y(n2050) );
  OAI21XL U1798 ( .A0(n982), .A1(n1706), .B0(n2051), .Y(n1300) );
  AOI2BB2X1 U1799 ( .B0(N1145), .B1(n1705), .A0N(n2015), .A1N(n985), .Y(n2051)
         );
  OAI221XL U1800 ( .A0(n979), .A1(n1698), .B0(n1531), .B1(n1697), .C0(n2052), 
        .Y(n1299) );
  AOI2BB2X1 U1801 ( .B0(n1696), .B1(\C1[3][1] ), .A0N(n1699), .A1N(n981), .Y(
        n2052) );
  OAI221XL U1802 ( .A0(n978), .A1(n1701), .B0(n1653), .B1(n1700), .C0(n2053), 
        .Y(n1298) );
  AOI2BB2X1 U1803 ( .B0(n2025), .B1(n1523), .A0N(n979), .A1N(n1702), .Y(n2053)
         );
  OAI222XL U1804 ( .A0(n1535), .A1(n1703), .B0(n979), .B1(n2028), .C0(n978), 
        .C1(n1704), .Y(n1297) );
  OAI221XL U1805 ( .A0(n977), .A1(n2007), .B0(n980), .B1(n1695), .C0(n2054), 
        .Y(n1296) );
  OAI21XL U1806 ( .A0(n977), .A1(n1706), .B0(n2055), .Y(n1295) );
  AOI2BB2X1 U1807 ( .B0(N1144), .B1(n1705), .A0N(n2015), .A1N(n980), .Y(n2055)
         );
  OAI21XL U1808 ( .A0(n1012), .A1(n1706), .B0(n2056), .Y(n1294) );
  AOI2BB2X1 U1809 ( .B0(N1150), .B1(n1705), .A0N(n2015), .A1N(n1013), .Y(n2056) );
  OAI221XL U1810 ( .A0(n2007), .A1(n1671), .B0(n1695), .B1(n1576), .C0(n2057), 
        .Y(n1293) );
  AOI22X1 U1811 ( .A0(n2612), .A1(n2010), .B0(n2011), .B1(\symbol[3][5] ), .Y(
        n2057) );
  OAI221XL U1812 ( .A0(n1698), .A1(n1504), .B0(n1479), .B1(n1697), .C0(n2058), 
        .Y(n1292) );
  OAI221XL U1813 ( .A0(n1701), .A1(n1558), .B0(n1487), .B1(n1700), .C0(n2060), 
        .Y(n1291) );
  AOI2BB2X1 U1814 ( .B0(n2612), .B1(n2025), .A0N(n1702), .A1N(n1504), .Y(n2060) );
  OAI222XL U1815 ( .A0(n1646), .A1(n1703), .B0(n2028), .B1(n1504), .C0(n1704), 
        .C1(n1558), .Y(n1290) );
  OAI222XL U1816 ( .A0(n2015), .A1(n1576), .B0(n2061), .B1(n2062), .C0(n1706), 
        .C1(n1671), .Y(n1289) );
  OAI221XL U1817 ( .A0(n2007), .A1(n1666), .B0(n1695), .B1(n1573), .C0(n2063), 
        .Y(n1288) );
  AOI22X1 U1818 ( .A0(n2613), .A1(n2010), .B0(n2011), .B1(\symbol[3][4] ), .Y(
        n2063) );
  OAI221XL U1819 ( .A0(n1698), .A1(n1505), .B0(n1483), .B1(n1697), .C0(n2064), 
        .Y(n1287) );
  OAI221XL U1820 ( .A0(n1701), .A1(n1559), .B0(n1516), .B1(n1700), .C0(n2065), 
        .Y(n1286) );
  AOI2BB2X1 U1821 ( .B0(n2613), .B1(n2025), .A0N(n1702), .A1N(n1505), .Y(n2065) );
  OAI222XL U1822 ( .A0(n1647), .A1(n1703), .B0(n2028), .B1(n1505), .C0(n1704), 
        .C1(n1559), .Y(n1285) );
  OAI221XL U1823 ( .A0(n2015), .A1(n1573), .B0(n1706), .B1(n1666), .C0(n2066), 
        .Y(n1284) );
  OAI21XL U1824 ( .A0(\symbol[4][4] ), .A1(\symbol[5][4] ), .B0(n1705), .Y(
        n2066) );
  OAI221XL U1825 ( .A0(n2007), .A1(n1667), .B0(n1695), .B1(n1574), .C0(n2067), 
        .Y(n1283) );
  AOI22X1 U1826 ( .A0(n2614), .A1(n2010), .B0(n2011), .B1(\symbol[3][3] ), .Y(
        n2067) );
  OAI221XL U1827 ( .A0(n1698), .A1(n1506), .B0(n1484), .B1(n1697), .C0(n2068), 
        .Y(n1282) );
  OAI221XL U1828 ( .A0(n1701), .A1(n1560), .B0(n1517), .B1(n1700), .C0(n2069), 
        .Y(n1281) );
  AOI2BB2X1 U1829 ( .B0(n2614), .B1(n2025), .A0N(n1702), .A1N(n1506), .Y(n2069) );
  OAI222XL U1830 ( .A0(n1648), .A1(n1703), .B0(n2028), .B1(n1506), .C0(n1704), 
        .C1(n1560), .Y(n1280) );
  OAI221XL U1831 ( .A0(n2015), .A1(n1574), .B0(n1706), .B1(n1667), .C0(n2070), 
        .Y(n1279) );
  OAI21XL U1832 ( .A0(\symbol[4][3] ), .A1(\symbol[5][3] ), .B0(n1705), .Y(
        n2070) );
  OAI221XL U1833 ( .A0(n2007), .A1(n1668), .B0(n1695), .B1(n1575), .C0(n2071), 
        .Y(n1278) );
  AOI22X1 U1834 ( .A0(n2615), .A1(n2010), .B0(n2011), .B1(\symbol[3][2] ), .Y(
        n2071) );
  OAI221XL U1835 ( .A0(n1698), .A1(n1507), .B0(n1485), .B1(n1697), .C0(n2072), 
        .Y(n1277) );
  OAI221XL U1836 ( .A0(n1701), .A1(n1561), .B0(n1518), .B1(n1700), .C0(n2073), 
        .Y(n1276) );
  AOI2BB2X1 U1837 ( .B0(n2615), .B1(n2025), .A0N(n1702), .A1N(n1507), .Y(n2073) );
  OAI222XL U1838 ( .A0(n1649), .A1(n1703), .B0(n2028), .B1(n1507), .C0(n1704), 
        .C1(n1561), .Y(n1275) );
  OAI221XL U1839 ( .A0(n2015), .A1(n1575), .B0(n1706), .B1(n1668), .C0(n2074), 
        .Y(n1274) );
  OAI21XL U1840 ( .A0(\symbol[4][2] ), .A1(\symbol[5][2] ), .B0(n1705), .Y(
        n2074) );
  OAI221XL U1841 ( .A0(n2007), .A1(n1669), .B0(n1695), .B1(n1571), .C0(n2075), 
        .Y(n1273) );
  AOI22X1 U1842 ( .A0(n2616), .A1(n2010), .B0(n2011), .B1(\symbol[3][1] ), .Y(
        n2075) );
  OAI221XL U1843 ( .A0(n1698), .A1(n1508), .B0(n1486), .B1(n1697), .C0(n2076), 
        .Y(n1272) );
  AOI22X1 U1844 ( .A0(n2610), .A1(n1696), .B0(n2616), .B1(n2059), .Y(n2076) );
  OAI221XL U1845 ( .A0(n1701), .A1(n1562), .B0(n1519), .B1(n1700), .C0(n2077), 
        .Y(n1271) );
  AOI2BB2X1 U1846 ( .B0(n2616), .B1(n2025), .A0N(n1702), .A1N(n1508), .Y(n2077) );
  OAI222XL U1847 ( .A0(n1650), .A1(n1703), .B0(n2028), .B1(n1508), .C0(n1704), 
        .C1(n1562), .Y(n1270) );
  OAI221XL U1848 ( .A0(n2015), .A1(n1571), .B0(n1706), .B1(n1669), .C0(n2078), 
        .Y(n1269) );
  OAI21XL U1849 ( .A0(\symbol[4][1] ), .A1(\symbol[5][1] ), .B0(n1705), .Y(
        n2078) );
  OAI221XL U1850 ( .A0(n2007), .A1(n1670), .B0(n1695), .B1(n1572), .C0(n2079), 
        .Y(n1268) );
  AOI22X1 U1851 ( .A0(n2617), .A1(n2010), .B0(n2011), .B1(\symbol[3][0] ), .Y(
        n2079) );
  OAI221XL U1852 ( .A0(n1698), .A1(n1509), .B0(n1482), .B1(n1697), .C0(n2082), 
        .Y(n1267) );
  AOI22X1 U1853 ( .A0(n2611), .A1(n1696), .B0(n2617), .B1(n2059), .Y(n2082) );
  CLKINVX1 U1854 ( .A(n1699), .Y(n2059) );
  OAI21XL U1855 ( .A0(n2080), .A1(n2083), .B0(n1825), .Y(n2085) );
  CLKINVX1 U1856 ( .A(n2081), .Y(n2080) );
  OAI22XL U1857 ( .A0(n1013), .A1(n1589), .B0(n2087), .B1(n2088), .Y(n2086) );
  NOR2X1 U1858 ( .A(n1011), .B(\C1[3][7] ), .Y(n2088) );
  AOI32X1 U1859 ( .A0(n2089), .A1(n2090), .A2(n2091), .B0(n2092), .B1(n2093), 
        .Y(n2087) );
  OAI21XL U1860 ( .A0(n2094), .A1(n1005), .B0(n1590), .Y(n2093) );
  NAND2X1 U1861 ( .A(n2094), .B(n1005), .Y(n2092) );
  AOI32X1 U1862 ( .A0(n996), .A1(\C1[3][4] ), .A2(n2090), .B0(\C1[3][5] ), 
        .B1(n1001), .Y(n2094) );
  AOI2BB2X1 U1863 ( .B0(n1525), .B1(n995), .A0N(\C1[3][6] ), .A1N(n1006), .Y(
        n2091) );
  NAND2X1 U1864 ( .A(n1000), .B(n1577), .Y(n2090) );
  OAI211X1 U1865 ( .A0(n990), .A1(n2095), .B0(n2096), .C0(n2097), .Y(n2089) );
  AO21X1 U1866 ( .A0(n2095), .A1(n990), .B0(n1524), .Y(n2097) );
  OAI222XL U1867 ( .A0(n991), .A1(\C1[3][3] ), .B0(n986), .B1(\C1[3][2] ), 
        .C0(n2098), .C1(n2099), .Y(n2096) );
  NAND2X1 U1868 ( .A(n986), .B(\C1[3][2] ), .Y(n2095) );
  OAI221XL U1869 ( .A0(n1701), .A1(n1563), .B0(n1520), .B1(n1700), .C0(n2100), 
        .Y(n1266) );
  AOI2BB2X1 U1870 ( .B0(n2617), .B1(n2025), .A0N(n1702), .A1N(n1509), .Y(n2100) );
  NOR2BX1 U1871 ( .AN(n2101), .B(n2102), .Y(n2083) );
  OAI22XL U1872 ( .A0(n1011), .A1(n1594), .B0(n2103), .B1(n2104), .Y(n2101) );
  NOR2X1 U1873 ( .A(n1010), .B(n1589), .Y(n2104) );
  AOI32X1 U1874 ( .A0(n2105), .A1(n2106), .A2(n2107), .B0(n2108), .B1(n2109), 
        .Y(n2103) );
  OAI21XL U1875 ( .A0(n2110), .A1(n1582), .B0(n1006), .Y(n2109) );
  NAND2X1 U1876 ( .A(n2110), .B(n1582), .Y(n2108) );
  AOI32X1 U1877 ( .A0(n994), .A1(n1525), .A2(n2106), .B0(n1577), .B1(n999), 
        .Y(n2110) );
  AOI2BB2X1 U1878 ( .B0(n996), .B1(n1526), .A0N(n1590), .A1N(n1004), .Y(n2107)
         );
  NAND2X1 U1879 ( .A(n1001), .B(n1584), .Y(n2106) );
  OAI211X1 U1880 ( .A0(n991), .A1(n2111), .B0(n2112), .C0(n2113), .Y(n2105) );
  AO21X1 U1881 ( .A0(n2111), .A1(n991), .B0(n1600), .Y(n2113) );
  OAI222XL U1882 ( .A0(n989), .A1(n1524), .B0(n984), .B1(n1578), .C0(n2114), 
        .C1(n2115), .Y(n2112) );
  CLKINVX1 U1883 ( .A(n2116), .Y(n2114) );
  NAND2X1 U1884 ( .A(n984), .B(n1578), .Y(n2111) );
  CLKINVX1 U1885 ( .A(n1822), .Y(n1825) );
  OAI222XL U1886 ( .A0(n1651), .A1(n1703), .B0(n2028), .B1(n1509), .C0(n1704), 
        .C1(n1563), .Y(n1265) );
  AOI2BB2X1 U1887 ( .B0(n1009), .B1(n1594), .A0N(n2118), .A1N(n2119), .Y(n2117) );
  NOR2X1 U1888 ( .A(n1009), .B(n1594), .Y(n2119) );
  AOI32X1 U1889 ( .A0(n2120), .A1(n2121), .A2(n2122), .B0(n2123), .B1(n2124), 
        .Y(n2118) );
  OAI21XL U1890 ( .A0(n2125), .A1(n1598), .B0(n1004), .Y(n2124) );
  NAND2X1 U1891 ( .A(n2125), .B(n1598), .Y(n2123) );
  AOI32X1 U1892 ( .A0(n993), .A1(n1526), .A2(n2121), .B0(n1584), .B1(n998), 
        .Y(n2125) );
  OA22X1 U1893 ( .A0(n1582), .A1(n1003), .B0(n1526), .B1(n993), .Y(n2122) );
  OR2X1 U1894 ( .A(n998), .B(n1584), .Y(n2121) );
  OAI211X1 U1895 ( .A0(n989), .A1(n2126), .B0(n2127), .C0(n2128), .Y(n2120) );
  OAI2BB1X1 U1896 ( .A0N(n2126), .A1N(n989), .B0(n988), .Y(n2128) );
  OAI222XL U1897 ( .A0(n988), .A1(n1600), .B0(n983), .B1(n1533), .C0(n2129), 
        .C1(n2130), .Y(n2127) );
  NOR2X1 U1898 ( .A(n979), .B(n1536), .Y(n2130) );
  AOI211X1 U1899 ( .A0(n979), .A1(n1536), .B0(n1602), .C0(n1008), .Y(n2129) );
  NAND2X1 U1900 ( .A(n983), .B(n1533), .Y(n2126) );
  CLKINVX1 U1901 ( .A(n1841), .Y(n1814) );
  NOR3X1 U1902 ( .A(n1581), .B(sort_stage[2]), .C(n1830), .Y(n1841) );
  OAI221XL U1903 ( .A0(n2015), .A1(n1572), .B0(n1706), .B1(n1670), .C0(n2131), 
        .Y(n1264) );
  OAI21XL U1904 ( .A0(\symbol[4][0] ), .A1(\symbol[5][0] ), .B0(n1705), .Y(
        n2131) );
  OA22X1 U1905 ( .A0(\C1[3][7] ), .A1(n1012), .B0(n2133), .B1(n2134), .Y(n2132) );
  NOR2BX1 U1906 ( .AN(n1012), .B(n1013), .Y(n2134) );
  AOI32X1 U1907 ( .A0(n2135), .A1(n2136), .A2(n2137), .B0(n2138), .B1(n2139), 
        .Y(n2133) );
  OAI21XL U1908 ( .A0(n2140), .A1(n1002), .B0(\C1[3][6] ), .Y(n2139) );
  NAND2X1 U1909 ( .A(n2140), .B(n1002), .Y(n2138) );
  AOI32X1 U1910 ( .A0(n995), .A1(\C1[4][4] ), .A2(n2136), .B0(\C1[4][5] ), 
        .B1(n1000), .Y(n2140) );
  AOI2BB2X1 U1911 ( .B0(\C1[3][6] ), .B1(n1002), .A0N(\C1[4][4] ), .A1N(n995), 
        .Y(n2137) );
  NAND2X1 U1912 ( .A(n997), .B(\C1[3][5] ), .Y(n2136) );
  OAI211X1 U1913 ( .A0(n987), .A1(n2141), .B0(n2142), .C0(n2143), .Y(n2135) );
  AO21X1 U1914 ( .A0(n2141), .A1(n987), .B0(\C1[3][3] ), .Y(n2143) );
  OAI222XL U1915 ( .A0(n990), .A1(\C1[4][3] ), .B0(n985), .B1(\C1[4][2] ), 
        .C0(n2144), .C1(n2145), .Y(n2142) );
  NOR2X1 U1916 ( .A(n977), .B(\C1[3][1] ), .Y(n2145) );
  AOI211X1 U1917 ( .A0(n977), .A1(\C1[3][1] ), .B0(\C1[3][0] ), .C0(n1015), 
        .Y(n2144) );
  NAND2X1 U1918 ( .A(n985), .B(\C1[4][2] ), .Y(n2141) );
  OAI221XL U1919 ( .A0(n944), .A1(n2146), .B0(n946), .B1(n1713), .C0(n2148), 
        .Y(n1263) );
  AOI2BB2X1 U1920 ( .B0(n2149), .B1(n1579), .A0N(n2150), .A1N(n945), .Y(n2148)
         );
  OAI21XL U1921 ( .A0(n945), .A1(n1714), .B0(n2152), .Y(n1262) );
  OAI221XL U1922 ( .A0(n941), .A1(n2146), .B0(n943), .B1(n1713), .C0(n2155), 
        .Y(n1261) );
  AOI2BB2X1 U1923 ( .B0(n2149), .B1(n1589), .A0N(n2150), .A1N(n942), .Y(n2155)
         );
  OAI221XL U1924 ( .A0(n940), .A1(n1716), .B0(n1010), .B1(n1715), .C0(n2158), 
        .Y(n1260) );
  AOI2BB2X1 U1925 ( .B0(n2159), .B1(\C2[2][7] ), .A0N(n941), .A1N(n1717), .Y(
        n2158) );
  OAI222XL U1926 ( .A0(n1009), .A1(n1718), .B0(n941), .B1(n2162), .C0(n940), 
        .C1(n1719), .Y(n1259) );
  OAI221XL U1927 ( .A0(n939), .A1(n1716), .B0(n1008), .B1(n1715), .C0(n2164), 
        .Y(n1258) );
  AOI2BB2X1 U1928 ( .B0(n2159), .B1(\C2[2][0] ), .A0N(n944), .A1N(n1717), .Y(
        n2164) );
  OAI221XL U1929 ( .A0(n936), .A1(n2146), .B0(n938), .B1(n1713), .C0(n2165), 
        .Y(n1257) );
  AOI2BB2X1 U1930 ( .B0(n2149), .B1(n1590), .A0N(n2150), .A1N(n937), .Y(n2165)
         );
  OAI221XL U1931 ( .A0(n935), .A1(n1716), .B0(n1004), .B1(n1715), .C0(n2166), 
        .Y(n1256) );
  AOI2BB2X1 U1932 ( .B0(n2159), .B1(\C2[2][6] ), .A0N(n936), .A1N(n1717), .Y(
        n2166) );
  OAI222XL U1933 ( .A0(n1003), .A1(n1718), .B0(n936), .B1(n2162), .C0(n935), 
        .C1(n1719), .Y(n1255) );
  OAI21XL U1934 ( .A0(n937), .A1(n1714), .B0(n2167), .Y(n1254) );
  OAI221XL U1935 ( .A0(n932), .A1(n2146), .B0(n934), .B1(n1713), .C0(n2168), 
        .Y(n1253) );
  AOI2BB2X1 U1936 ( .B0(n2149), .B1(n1577), .A0N(n2150), .A1N(n933), .Y(n2168)
         );
  OAI221XL U1937 ( .A0(n931), .A1(n1716), .B0(n999), .B1(n1715), .C0(n2169), 
        .Y(n1252) );
  AOI2BB2X1 U1938 ( .B0(n2159), .B1(\C2[2][5] ), .A0N(n932), .A1N(n1717), .Y(
        n2169) );
  OAI222XL U1939 ( .A0(n998), .A1(n1718), .B0(n932), .B1(n2162), .C0(n931), 
        .C1(n1719), .Y(n1251) );
  OAI21XL U1940 ( .A0(n933), .A1(n1714), .B0(n2170), .Y(n1250) );
  OAI221XL U1941 ( .A0(n928), .A1(n2146), .B0(n930), .B1(n1713), .C0(n2171), 
        .Y(n1249) );
  AOI2BB2X1 U1942 ( .B0(n2149), .B1(n1525), .A0N(n2150), .A1N(n929), .Y(n2171)
         );
  OAI221XL U1943 ( .A0(n927), .A1(n1716), .B0(n994), .B1(n1715), .C0(n2172), 
        .Y(n1248) );
  AOI2BB2X1 U1944 ( .B0(n2159), .B1(\C2[2][4] ), .A0N(n928), .A1N(n1717), .Y(
        n2172) );
  OAI222XL U1945 ( .A0(n993), .A1(n1718), .B0(n928), .B1(n2162), .C0(n927), 
        .C1(n1719), .Y(n1247) );
  OAI21XL U1946 ( .A0(n929), .A1(n1714), .B0(n2173), .Y(n1246) );
  OAI221XL U1947 ( .A0(n924), .A1(n2146), .B0(n926), .B1(n1713), .C0(n2174), 
        .Y(n1245) );
  AOI2BB2X1 U1948 ( .B0(n2149), .B1(n1524), .A0N(n2150), .A1N(n925), .Y(n2174)
         );
  OAI221XL U1949 ( .A0(n923), .A1(n1716), .B0(n989), .B1(n1715), .C0(n2175), 
        .Y(n1244) );
  AOI2BB2X1 U1950 ( .B0(n2159), .B1(\C2[2][3] ), .A0N(n924), .A1N(n1717), .Y(
        n2175) );
  OAI222XL U1951 ( .A0(n988), .A1(n1718), .B0(n924), .B1(n2162), .C0(n923), 
        .C1(n1719), .Y(n1243) );
  OAI21XL U1952 ( .A0(n925), .A1(n1714), .B0(n2176), .Y(n1242) );
  OAI221XL U1953 ( .A0(n920), .A1(n2146), .B0(n922), .B1(n1713), .C0(n2177), 
        .Y(n1241) );
  AOI2BB2X1 U1954 ( .B0(n2149), .B1(n1578), .A0N(n2150), .A1N(n921), .Y(n2177)
         );
  OAI221XL U1955 ( .A0(n919), .A1(n1716), .B0(n984), .B1(n1715), .C0(n2178), 
        .Y(n1240) );
  AOI2BB2X1 U1956 ( .B0(n2159), .B1(\C2[2][2] ), .A0N(n920), .A1N(n1717), .Y(
        n2178) );
  OAI222XL U1957 ( .A0(n983), .A1(n1718), .B0(n920), .B1(n2162), .C0(n919), 
        .C1(n1719), .Y(n1239) );
  OAI21XL U1958 ( .A0(n921), .A1(n1714), .B0(n2179), .Y(n1238) );
  OAI221XL U1959 ( .A0(n916), .A1(n2146), .B0(n918), .B1(n1713), .C0(n2180), 
        .Y(n1237) );
  AOI2BB2X1 U1960 ( .B0(n2149), .B1(n1523), .A0N(n2150), .A1N(n917), .Y(n2180)
         );
  OAI221XL U1961 ( .A0(n915), .A1(n1716), .B0(n979), .B1(n1715), .C0(n2181), 
        .Y(n1236) );
  AOI2BB2X1 U1962 ( .B0(n2159), .B1(\C2[2][1] ), .A0N(n916), .A1N(n1717), .Y(
        n2181) );
  OAI222XL U1963 ( .A0(n978), .A1(n1718), .B0(n916), .B1(n2162), .C0(n915), 
        .C1(n1719), .Y(n1235) );
  OAI21XL U1964 ( .A0(n917), .A1(n1714), .B0(n2182), .Y(n1234) );
  OAI222XL U1965 ( .A0(n1007), .A1(n1718), .B0(n944), .B1(n2162), .C0(n939), 
        .C1(n1719), .Y(n1233) );
  OAI21XL U1966 ( .A0(n942), .A1(n1714), .B0(n2183), .Y(n1232) );
  OAI222XL U1967 ( .A0(n1721), .A1(n914), .B0(n2186), .B1(n1720), .C0(n2188), 
        .C1(n913), .Y(n1231) );
  CLKINVX1 U1968 ( .A(N2261), .Y(n2186) );
  OAI221XL U1969 ( .A0(n914), .A1(n2189), .B0(n941), .B1(n1723), .C0(n2191), 
        .Y(n1230) );
  OA22X1 U1970 ( .A0(n912), .A1(n1722), .B0(n913), .B1(n1724), .Y(n2191) );
  OAI222XL U1971 ( .A0(n940), .A1(n1725), .B0(n913), .B1(n2195), .C0(n912), 
        .C1(n1726), .Y(n1229) );
  OAI221XL U1972 ( .A0(n910), .A1(n2189), .B0(n944), .B1(n1723), .C0(n2197), 
        .Y(n1228) );
  OA22X1 U1973 ( .A0(n909), .A1(n1722), .B0(n911), .B1(n1724), .Y(n2197) );
  OAI222XL U1974 ( .A0(n939), .A1(n1725), .B0(n911), .B1(n2195), .C0(n909), 
        .C1(n1726), .Y(n1227) );
  OAI222XL U1975 ( .A0(n1721), .A1(n910), .B0(n2198), .B1(n1720), .C0(n2188), 
        .C1(n911), .Y(n1226) );
  CLKINVX1 U1976 ( .A(N2254), .Y(n2198) );
  OAI222XL U1977 ( .A0(n1721), .A1(n908), .B0(n2199), .B1(n1720), .C0(n2188), 
        .C1(n907), .Y(n1225) );
  CLKINVX1 U1978 ( .A(N2255), .Y(n2199) );
  OAI221XL U1979 ( .A0(n908), .A1(n2189), .B0(n916), .B1(n1723), .C0(n2200), 
        .Y(n1224) );
  OA22X1 U1980 ( .A0(n906), .A1(n1722), .B0(n907), .B1(n1724), .Y(n2200) );
  OAI222XL U1981 ( .A0(n915), .A1(n1725), .B0(n907), .B1(n2195), .C0(n906), 
        .C1(n1726), .Y(n1223) );
  OAI222XL U1982 ( .A0(n1721), .A1(n905), .B0(n2201), .B1(n1720), .C0(n2188), 
        .C1(n904), .Y(n1222) );
  CLKINVX1 U1983 ( .A(N2256), .Y(n2201) );
  OAI221XL U1984 ( .A0(n905), .A1(n2189), .B0(n920), .B1(n1723), .C0(n2202), 
        .Y(n1221) );
  OA22X1 U1985 ( .A0(n903), .A1(n1722), .B0(n904), .B1(n1724), .Y(n2202) );
  OAI222XL U1986 ( .A0(n919), .A1(n1725), .B0(n904), .B1(n2195), .C0(n903), 
        .C1(n1726), .Y(n1220) );
  OAI222XL U1987 ( .A0(n1721), .A1(n902), .B0(n2203), .B1(n1720), .C0(n2188), 
        .C1(n901), .Y(n1219) );
  CLKINVX1 U1988 ( .A(N2257), .Y(n2203) );
  OAI221XL U1989 ( .A0(n902), .A1(n2189), .B0(n924), .B1(n1723), .C0(n2204), 
        .Y(n1218) );
  OA22X1 U1990 ( .A0(n900), .A1(n1722), .B0(n901), .B1(n1724), .Y(n2204) );
  OAI222XL U1991 ( .A0(n923), .A1(n1725), .B0(n901), .B1(n2195), .C0(n900), 
        .C1(n1726), .Y(n1217) );
  OAI222XL U1992 ( .A0(n1721), .A1(n899), .B0(n2205), .B1(n1720), .C0(n2188), 
        .C1(n898), .Y(n1216) );
  CLKINVX1 U1993 ( .A(N2258), .Y(n2205) );
  OAI221XL U1994 ( .A0(n899), .A1(n2189), .B0(n928), .B1(n1723), .C0(n2206), 
        .Y(n1215) );
  OA22X1 U1995 ( .A0(n897), .A1(n1722), .B0(n898), .B1(n1724), .Y(n2206) );
  OAI222XL U1996 ( .A0(n927), .A1(n1725), .B0(n898), .B1(n2195), .C0(n897), 
        .C1(n1726), .Y(n1214) );
  OAI222XL U1997 ( .A0(n1721), .A1(n896), .B0(n2207), .B1(n1720), .C0(n2188), 
        .C1(n895), .Y(n1213) );
  CLKINVX1 U1998 ( .A(N2259), .Y(n2207) );
  OAI221XL U1999 ( .A0(n896), .A1(n2189), .B0(n932), .B1(n1723), .C0(n2208), 
        .Y(n1212) );
  OA22X1 U2000 ( .A0(n894), .A1(n1722), .B0(n895), .B1(n1724), .Y(n2208) );
  OAI222XL U2001 ( .A0(n931), .A1(n1725), .B0(n895), .B1(n2195), .C0(n894), 
        .C1(n1726), .Y(n1211) );
  OAI222XL U2002 ( .A0(n1721), .A1(n893), .B0(n2209), .B1(n1720), .C0(n2188), 
        .C1(n892), .Y(n1210) );
  CLKINVX1 U2003 ( .A(N2260), .Y(n2209) );
  OAI221XL U2004 ( .A0(n893), .A1(n2189), .B0(n936), .B1(n1723), .C0(n2210), 
        .Y(n1209) );
  OA22X1 U2005 ( .A0(n891), .A1(n1722), .B0(n892), .B1(n1724), .Y(n2210) );
  OAI222XL U2006 ( .A0(n935), .A1(n1725), .B0(n892), .B1(n2195), .C0(n891), 
        .C1(n1726), .Y(n1208) );
  OAI222XL U2007 ( .A0(n912), .A1(n1735), .B0(n889), .B1(n1738), .C0(n890), 
        .C1(n1740), .Y(n1207) );
  OAI222XL U2008 ( .A0(n1736), .A1(n2212), .B0(n890), .B1(n1738), .C0(n889), 
        .C1(n1740), .Y(n1206) );
  CLKINVX1 U2009 ( .A(N2782), .Y(n2212) );
  OAI222XL U2010 ( .A0(n909), .A1(n1735), .B0(n887), .B1(n1738), .C0(n888), 
        .C1(n1740), .Y(n1205) );
  OAI222XL U2011 ( .A0(n1736), .A1(n2213), .B0(n888), .B1(n1738), .C0(n887), 
        .C1(n1740), .Y(n1204) );
  CLKINVX1 U2012 ( .A(N2775), .Y(n2213) );
  OAI222XL U2013 ( .A0(n906), .A1(n1735), .B0(n885), .B1(n1738), .C0(n886), 
        .C1(n1740), .Y(n1203) );
  OAI222XL U2014 ( .A0(n1736), .A1(n2214), .B0(n886), .B1(n1738), .C0(n885), 
        .C1(n1740), .Y(n1202) );
  CLKINVX1 U2015 ( .A(N2776), .Y(n2214) );
  OAI222XL U2016 ( .A0(n903), .A1(n1735), .B0(n883), .B1(n1738), .C0(n884), 
        .C1(n1740), .Y(n1201) );
  OAI222XL U2017 ( .A0(n1736), .A1(n2215), .B0(n884), .B1(n1738), .C0(n883), 
        .C1(n1740), .Y(n1200) );
  CLKINVX1 U2018 ( .A(N2777), .Y(n2215) );
  OAI222XL U2019 ( .A0(n900), .A1(n1735), .B0(n881), .B1(n1738), .C0(n882), 
        .C1(n1740), .Y(n1199) );
  OAI222XL U2020 ( .A0(n1736), .A1(n2216), .B0(n882), .B1(n1738), .C0(n881), 
        .C1(n1740), .Y(n1198) );
  CLKINVX1 U2021 ( .A(N2778), .Y(n2216) );
  OAI222XL U2022 ( .A0(n897), .A1(n1735), .B0(n879), .B1(n1738), .C0(n880), 
        .C1(n1740), .Y(n1197) );
  OAI222XL U2023 ( .A0(n1736), .A1(n2217), .B0(n880), .B1(n1738), .C0(n879), 
        .C1(n1740), .Y(n1196) );
  CLKINVX1 U2024 ( .A(N2779), .Y(n2217) );
  OAI222XL U2025 ( .A0(n894), .A1(n1735), .B0(n877), .B1(n1738), .C0(n878), 
        .C1(n1740), .Y(n1195) );
  OAI222XL U2026 ( .A0(n1736), .A1(n2218), .B0(n878), .B1(n1480), .C0(n877), 
        .C1(n1740), .Y(n1194) );
  CLKINVX1 U2027 ( .A(N2780), .Y(n2218) );
  OAI222XL U2028 ( .A0(n891), .A1(n1735), .B0(n875), .B1(n1738), .C0(n876), 
        .C1(n1740), .Y(n1193) );
  OAI222XL U2029 ( .A0(n1736), .A1(n2219), .B0(n876), .B1(n1737), .C0(n875), 
        .C1(n1740), .Y(n1192) );
  CLKINVX1 U2030 ( .A(N2781), .Y(n2219) );
  OAI222XL U2031 ( .A0(n2154), .A1(n1660), .B0(n2220), .B1(n2184), .C0(n1714), 
        .C1(n1546), .Y(n1191) );
  OAI221XL U2032 ( .A0(n2146), .A1(n1510), .B0(n1713), .B1(n1660), .C0(n2221), 
        .Y(n1190) );
  AOI2BB2X1 U2033 ( .B0(n2149), .B1(n2612), .A0N(n1546), .A1N(n2150), .Y(n2221) );
  OAI221XL U2034 ( .A0(n1716), .A1(n1640), .B0(n1504), .B1(n1715), .C0(n2222), 
        .Y(n1189) );
  AOI2BB2X1 U2035 ( .B0(n2593), .B1(n2159), .A0N(n1717), .A1N(n1510), .Y(n2222) );
  OAI222XL U2036 ( .A0(n1558), .A1(n1718), .B0(n2162), .B1(n1510), .C0(n1719), 
        .C1(n1640), .Y(n1188) );
  OAI222XL U2037 ( .A0(n2188), .A1(n1497), .B0(n2223), .B1(n1720), .C0(n1721), 
        .C1(n1672), .Y(n1187) );
  OAI221XL U2038 ( .A0(n2189), .A1(n1672), .B0(n1723), .B1(n1510), .C0(n2224), 
        .Y(n1186) );
  OA22X1 U2039 ( .A0(n1722), .A1(n1565), .B0(n1724), .B1(n1497), .Y(n2224) );
  OAI222XL U2040 ( .A0(n1725), .A1(n1640), .B0(n2195), .B1(n1497), .C0(n1726), 
        .C1(n1565), .Y(n1185) );
  OAI222XL U2041 ( .A0(n1737), .A1(n1678), .B0(n2225), .B1(n1735), .C0(n1740), 
        .C1(n1503), .Y(n1184) );
  OAI222XL U2042 ( .A0(n1736), .A1(n1565), .B0(n1737), .B1(n1503), .C0(n1739), 
        .C1(n1678), .Y(n1183) );
  XNOR2X1 U2043 ( .A(n2513), .B(n2226), .Y(n1182) );
  XNOR2X1 U2044 ( .A(n1637), .B(n2227), .Y(n1180) );
  NOR2X1 U2045 ( .A(n2226), .B(n2228), .Y(n2227) );
  OAI22XL U2046 ( .A0(n2228), .A1(n2229), .B0(n2509), .B1(n2230), .Y(n1179) );
  OA21XL U2047 ( .A0(n1708), .A1(n2232), .B0(n2233), .Y(n2230) );
  OAI22XL U2048 ( .A0(n2229), .A1(n1804), .B0(n2510), .B1(n2234), .Y(n1178) );
  OA21XL U2049 ( .A0(n1708), .A1(n2235), .B0(n2233), .Y(n2234) );
  OAI22XL U2050 ( .A0(n2236), .A1(n2229), .B0(n2512), .B1(n2237), .Y(n1177) );
  OA21XL U2051 ( .A0(n1708), .A1(n1805), .B0(n2233), .Y(n2237) );
  OAI22XL U2052 ( .A0(n2229), .A1(n2238), .B0(n2514), .B1(n2239), .Y(n1176) );
  OA21XL U2053 ( .A0(n1708), .A1(n2240), .B0(n2233), .Y(n2239) );
  NAND2X1 U2054 ( .A(n2241), .B(n1637), .Y(n2229) );
  OAI22XL U2055 ( .A0(n2228), .A1(n2242), .B0(n2505), .B1(n2243), .Y(n1175) );
  OA21XL U2056 ( .A0(n1708), .A1(n2232), .B0(n2244), .Y(n2243) );
  CLKINVX1 U2057 ( .A(n2232), .Y(n2228) );
  NOR2X1 U2058 ( .A(n1552), .B(n1638), .Y(n2232) );
  OAI22XL U2059 ( .A0(n1804), .A1(n2242), .B0(n2506), .B1(n2245), .Y(n1174) );
  OA21XL U2060 ( .A0(n1708), .A1(n2235), .B0(n2244), .Y(n2245) );
  CLKINVX1 U2061 ( .A(n2235), .Y(n1804) );
  NOR2X1 U2062 ( .A(n1638), .B(n2513), .Y(n2235) );
  OAI22XL U2063 ( .A0(n2236), .A1(n2242), .B0(n2507), .B1(n2246), .Y(n1173) );
  OA21XL U2064 ( .A0(n1708), .A1(n1805), .B0(n2244), .Y(n2246) );
  CLKINVX1 U2065 ( .A(n1805), .Y(n2236) );
  NOR2X1 U2066 ( .A(n1552), .B(n2511), .Y(n1805) );
  OAI22XL U2067 ( .A0(n2238), .A1(n2242), .B0(n2508), .B1(n2247), .Y(n1172) );
  OA21XL U2068 ( .A0(n1708), .A1(n2240), .B0(n2244), .Y(n2247) );
  NAND2X1 U2069 ( .A(n2515), .B(n2241), .Y(n2242) );
  AO22X1 U2070 ( .A0(n2248), .A1(n2249), .B0(n2250), .B1(n1707), .Y(n2241) );
  OAI22XL U2071 ( .A0(n1730), .A1(n1503), .B0(n1729), .B1(n1546), .Y(n2250) );
  OAI22XL U2072 ( .A0(n2606), .A1(n1728), .B0(n2580), .B1(n1828), .Y(n2248) );
  CLKINVX1 U2073 ( .A(n2240), .Y(n2238) );
  NOR2X1 U2074 ( .A(n2513), .B(n2511), .Y(n2240) );
  NAND2X1 U2075 ( .A(n862), .B(n2226), .Y(n1171) );
  OAI22XL U2076 ( .A0(n861), .A1(n1707), .B0(n862), .B1(n2251), .Y(n1170) );
  OAI22XL U2077 ( .A0(n860), .A1(n1707), .B0(n861), .B1(n2251), .Y(n1169) );
  OAI22XL U2078 ( .A0(n859), .A1(n1707), .B0(n860), .B1(n2251), .Y(n1168) );
  OAI22XL U2079 ( .A0(n858), .A1(n1707), .B0(n859), .B1(n2251), .Y(n1167) );
  OAI22XL U2080 ( .A0(n857), .A1(n1707), .B0(n858), .B1(n2251), .Y(n1166) );
  OAI22XL U2081 ( .A0(n856), .A1(n1707), .B0(n857), .B1(n2251), .Y(n1165) );
  OAI22XL U2082 ( .A0(n855), .A1(n1707), .B0(n856), .B1(n2251), .Y(n1164) );
  NAND2X1 U2083 ( .A(n2252), .B(n1707), .Y(n2251) );
  NOR2X1 U2084 ( .A(n2249), .B(n1708), .Y(n2226) );
  NOR2X1 U2085 ( .A(\symbol[5][5] ), .B(\symbol[4][5] ), .Y(n2061) );
  NOR2X1 U2086 ( .A(n2600), .B(n2606), .Y(n2220) );
  NOR2X1 U2087 ( .A(n2587), .B(n2593), .Y(n2223) );
  OAI21XL U2088 ( .A0(n2562), .A1(n2561), .B0(n2259), .Y(n2255) );
  NOR2X1 U2089 ( .A(n2574), .B(n2580), .Y(n2225) );
  OAI222XL U2090 ( .A0(n2154), .A1(n1661), .B0(n2260), .B1(n2184), .C0(n1714), 
        .C1(n1547), .Y(n1163) );
  OAI221XL U2091 ( .A0(n2146), .A1(n1511), .B0(n1713), .B1(n1661), .C0(n2261), 
        .Y(n1162) );
  AOI2BB2X1 U2092 ( .B0(n2149), .B1(n2613), .A0N(n1547), .A1N(n2150), .Y(n2261) );
  OAI221XL U2093 ( .A0(n1716), .A1(n1641), .B0(n1505), .B1(n1715), .C0(n2262), 
        .Y(n1161) );
  AOI2BB2X1 U2094 ( .B0(n2594), .B1(n2159), .A0N(n1717), .A1N(n1511), .Y(n2262) );
  OAI222XL U2095 ( .A0(n1559), .A1(n1718), .B0(n2162), .B1(n1511), .C0(n1719), 
        .C1(n1641), .Y(n1160) );
  OAI222XL U2096 ( .A0(n2188), .A1(n1498), .B0(n2263), .B1(n1720), .C0(n1721), 
        .C1(n1673), .Y(n1159) );
  OAI221XL U2097 ( .A0(n2189), .A1(n1673), .B0(n1723), .B1(n1511), .C0(n2264), 
        .Y(n1158) );
  OA22X1 U2098 ( .A0(n1722), .A1(n1566), .B0(n1724), .B1(n1498), .Y(n2264) );
  OAI222XL U2099 ( .A0(n1725), .A1(n1641), .B0(n2195), .B1(n1498), .C0(n1726), 
        .C1(n1566), .Y(n1157) );
  OAI222XL U2100 ( .A0(n1737), .A1(n1679), .B0(n2265), .B1(n1735), .C0(n1739), 
        .C1(n1488), .Y(n1156) );
  OAI222XL U2101 ( .A0(n1736), .A1(n1566), .B0(n1737), .B1(n1488), .C0(n1739), 
        .C1(n1679), .Y(n1155) );
  XNOR2X1 U2102 ( .A(n2523), .B(n2266), .Y(n1154) );
  XNOR2X1 U2103 ( .A(n1632), .B(n2267), .Y(n1152) );
  NOR2X1 U2104 ( .A(n2266), .B(n2268), .Y(n2267) );
  OAI22XL U2105 ( .A0(n2268), .A1(n2269), .B0(n2519), .B1(n2270), .Y(n1151) );
  OAI22XL U2106 ( .A0(n2269), .A1(n1800), .B0(n2520), .B1(n2273), .Y(n1150) );
  OAI22XL U2107 ( .A0(n2274), .A1(n2269), .B0(n2522), .B1(n2275), .Y(n1149) );
  OR3X1 U2108 ( .A(n2269), .B(n2523), .C(n2521), .Y(n2278) );
  NAND2X1 U2109 ( .A(n2279), .B(n1632), .Y(n2269) );
  OAI21XL U2110 ( .A0(n2280), .A1(n2272), .B0(HC5[0]), .Y(n2277) );
  OAI22XL U2111 ( .A0(n2268), .A1(n2281), .B0(n2516), .B1(n2282), .Y(n1147) );
  NAND2X1 U2112 ( .A(n2523), .B(n2521), .Y(n2268) );
  OAI22XL U2113 ( .A0(n1800), .A1(n2281), .B0(n2517), .B1(n2284), .Y(n1146) );
  NAND2X1 U2114 ( .A(n2521), .B(n1627), .Y(n1800) );
  OAI22XL U2115 ( .A0(n2274), .A1(n2281), .B0(n2518), .B1(n2285), .Y(n1145) );
  CLKINVX1 U2116 ( .A(n1801), .Y(n2274) );
  NOR2X1 U2117 ( .A(n1627), .B(n2521), .Y(n1801) );
  OAI31XL U2118 ( .A0(n2281), .A1(n2521), .A2(n2523), .B0(n2286), .Y(n1144) );
  OAI21XL U2119 ( .A0(n2280), .A1(n2283), .B0(HC5[4]), .Y(n2286) );
  OA21XL U2120 ( .A0(n2523), .A1(n2521), .B0(n2271), .Y(n2280) );
  NAND2X1 U2121 ( .A(n2524), .B(n2279), .Y(n2281) );
  AO22X1 U2122 ( .A0(n2287), .A1(n2288), .B0(n2289), .B1(n1709), .Y(n2279) );
  OAI22XL U2123 ( .A0(n1730), .A1(n1488), .B0(n1729), .B1(n1547), .Y(n2289) );
  OAI22XL U2124 ( .A0(n2607), .A1(n1728), .B0(n2581), .B1(n1828), .Y(n2287) );
  NAND2X1 U2125 ( .A(n841), .B(n2266), .Y(n1143) );
  OAI22XL U2126 ( .A0(n840), .A1(n1709), .B0(n841), .B1(n2290), .Y(n1142) );
  OAI22XL U2127 ( .A0(n839), .A1(n1709), .B0(n840), .B1(n2290), .Y(n1141) );
  OAI22XL U2128 ( .A0(n838), .A1(n1709), .B0(n839), .B1(n2290), .Y(n1140) );
  OAI22XL U2129 ( .A0(n837), .A1(n1709), .B0(n838), .B1(n2290), .Y(n1139) );
  OAI22XL U2130 ( .A0(n836), .A1(n1709), .B0(n837), .B1(n2290), .Y(n1138) );
  OAI22XL U2131 ( .A0(n835), .A1(n1709), .B0(n836), .B1(n2290), .Y(n1137) );
  OAI22XL U2132 ( .A0(n834), .A1(n1709), .B0(n835), .B1(n2290), .Y(n1136) );
  NAND2X1 U2133 ( .A(n2252), .B(n1709), .Y(n2290) );
  NOR2X1 U2134 ( .A(n2288), .B(n2276), .Y(n2266) );
  NOR2X1 U2135 ( .A(n2601), .B(n2607), .Y(n2260) );
  NOR2X1 U2136 ( .A(n2588), .B(n2594), .Y(n2263) );
  OAI21XL U2137 ( .A0(n2564), .A1(n2563), .B0(n2259), .Y(n2291) );
  NOR2X1 U2138 ( .A(n2575), .B(n2581), .Y(n2265) );
  OAI222XL U2139 ( .A0(n2154), .A1(n1662), .B0(n2293), .B1(n2184), .C0(n1714), 
        .C1(n1548), .Y(n1135) );
  OAI221XL U2140 ( .A0(n2146), .A1(n1512), .B0(n1713), .B1(n1662), .C0(n2294), 
        .Y(n1134) );
  AOI2BB2X1 U2141 ( .B0(n2149), .B1(n2614), .A0N(n1548), .A1N(n2150), .Y(n2294) );
  OAI221XL U2142 ( .A0(n1716), .A1(n1642), .B0(n1506), .B1(n1715), .C0(n2295), 
        .Y(n1133) );
  AOI2BB2X1 U2143 ( .B0(n2595), .B1(n2159), .A0N(n1717), .A1N(n1512), .Y(n2295) );
  OAI222XL U2144 ( .A0(n1560), .A1(n1718), .B0(n2162), .B1(n1512), .C0(n1719), 
        .C1(n1642), .Y(n1132) );
  OAI222XL U2145 ( .A0(n2188), .A1(n1499), .B0(n2296), .B1(n1720), .C0(n1721), 
        .C1(n1674), .Y(n1131) );
  OAI221XL U2146 ( .A0(n2189), .A1(n1674), .B0(n1723), .B1(n1512), .C0(n2297), 
        .Y(n1130) );
  OA22X1 U2147 ( .A0(n1722), .A1(n1567), .B0(n1724), .B1(n1499), .Y(n2297) );
  OAI222XL U2148 ( .A0(n1725), .A1(n1642), .B0(n2195), .B1(n1499), .C0(n1726), 
        .C1(n1567), .Y(n1129) );
  OAI222XL U2149 ( .A0(n1737), .A1(n1680), .B0(n2298), .B1(n1735), .C0(n1739), 
        .C1(n1489), .Y(n1128) );
  OAI222XL U2150 ( .A0(n1735), .A1(n1567), .B0(n1737), .B1(n1489), .C0(n1739), 
        .C1(n1680), .Y(n1127) );
  XNOR2X1 U2151 ( .A(n2532), .B(n2299), .Y(n1126) );
  XNOR2X1 U2152 ( .A(n1633), .B(n2300), .Y(n1124) );
  NOR2X1 U2153 ( .A(n2299), .B(n2301), .Y(n2300) );
  OAI22XL U2154 ( .A0(n2301), .A1(n2302), .B0(n2528), .B1(n2303), .Y(n1123) );
  OAI22XL U2155 ( .A0(n2302), .A1(n1796), .B0(n2529), .B1(n2306), .Y(n1122) );
  OAI22XL U2156 ( .A0(n2307), .A1(n2302), .B0(n2531), .B1(n2308), .Y(n1121) );
  OR3X1 U2157 ( .A(n2302), .B(n2532), .C(n2530), .Y(n2311) );
  NAND2X1 U2158 ( .A(n2312), .B(n1633), .Y(n2302) );
  OAI21XL U2159 ( .A0(n2313), .A1(n2305), .B0(HC4[0]), .Y(n2310) );
  OAI22XL U2160 ( .A0(n2301), .A1(n2314), .B0(n2525), .B1(n2315), .Y(n1119) );
  NAND2X1 U2161 ( .A(n2532), .B(n2530), .Y(n2301) );
  OAI22XL U2162 ( .A0(n1796), .A1(n2314), .B0(n2526), .B1(n2317), .Y(n1118) );
  NAND2X1 U2163 ( .A(n2530), .B(n1628), .Y(n1796) );
  OAI22XL U2164 ( .A0(n2307), .A1(n2314), .B0(n2527), .B1(n2318), .Y(n1117) );
  CLKINVX1 U2165 ( .A(n1797), .Y(n2307) );
  NOR2X1 U2166 ( .A(n1628), .B(n2530), .Y(n1797) );
  OAI31XL U2167 ( .A0(n2314), .A1(n2530), .A2(n2532), .B0(n2319), .Y(n1116) );
  OAI21XL U2168 ( .A0(n2313), .A1(n2316), .B0(HC4[4]), .Y(n2319) );
  OA21XL U2169 ( .A0(n2532), .A1(n2530), .B0(n2304), .Y(n2313) );
  NAND2X1 U2170 ( .A(n2533), .B(n2312), .Y(n2314) );
  AO22X1 U2171 ( .A0(n2320), .A1(n2321), .B0(n2322), .B1(n1710), .Y(n2312) );
  OAI22XL U2172 ( .A0(n1730), .A1(n1489), .B0(n1729), .B1(n1548), .Y(n2322) );
  OAI22XL U2173 ( .A0(n2608), .A1(n1728), .B0(n2582), .B1(n1828), .Y(n2320) );
  NAND2X1 U2174 ( .A(n820), .B(n2299), .Y(n1115) );
  OAI22XL U2175 ( .A0(n819), .A1(n1710), .B0(n820), .B1(n2323), .Y(n1114) );
  OAI22XL U2176 ( .A0(n818), .A1(n1710), .B0(n819), .B1(n2323), .Y(n1113) );
  OAI22XL U2177 ( .A0(n817), .A1(n1710), .B0(n818), .B1(n2323), .Y(n1112) );
  OAI22XL U2178 ( .A0(n816), .A1(n1710), .B0(n817), .B1(n2323), .Y(n1111) );
  OAI22XL U2179 ( .A0(n815), .A1(n1710), .B0(n816), .B1(n2323), .Y(n1110) );
  OAI22XL U2180 ( .A0(n814), .A1(n1710), .B0(n815), .B1(n2323), .Y(n1109) );
  OAI22XL U2181 ( .A0(n813), .A1(n1710), .B0(n814), .B1(n2323), .Y(n1108) );
  NAND2X1 U2182 ( .A(n2252), .B(n1710), .Y(n2323) );
  NOR2X1 U2183 ( .A(n2321), .B(n2309), .Y(n2299) );
  NOR2X1 U2184 ( .A(n2602), .B(n2608), .Y(n2293) );
  NOR2X1 U2185 ( .A(n2589), .B(n2595), .Y(n2296) );
  OAI21XL U2186 ( .A0(n2566), .A1(n2565), .B0(n2259), .Y(n2324) );
  NOR2X1 U2187 ( .A(n2576), .B(n2582), .Y(n2298) );
  OAI222XL U2188 ( .A0(n2154), .A1(n1663), .B0(n2326), .B1(n2184), .C0(n1714), 
        .C1(n1549), .Y(n1107) );
  OAI221XL U2189 ( .A0(n2146), .A1(n1513), .B0(n1713), .B1(n1663), .C0(n2327), 
        .Y(n1106) );
  AOI2BB2X1 U2190 ( .B0(n2149), .B1(n2615), .A0N(n1549), .A1N(n2150), .Y(n2327) );
  OAI221XL U2191 ( .A0(n1716), .A1(n1643), .B0(n1507), .B1(n1715), .C0(n2328), 
        .Y(n1105) );
  AOI2BB2X1 U2192 ( .B0(n2596), .B1(n2159), .A0N(n1717), .A1N(n1513), .Y(n2328) );
  OAI222XL U2193 ( .A0(n1561), .A1(n1718), .B0(n2162), .B1(n1513), .C0(n1719), 
        .C1(n1643), .Y(n1104) );
  OAI222XL U2194 ( .A0(n2188), .A1(n1500), .B0(n2329), .B1(n1720), .C0(n1721), 
        .C1(n1675), .Y(n1103) );
  OAI221XL U2195 ( .A0(n2189), .A1(n1675), .B0(n1723), .B1(n1513), .C0(n2330), 
        .Y(n1102) );
  OA22X1 U2196 ( .A0(n1722), .A1(n1568), .B0(n1724), .B1(n1500), .Y(n2330) );
  OAI222XL U2197 ( .A0(n1725), .A1(n1643), .B0(n2195), .B1(n1500), .C0(n1726), 
        .C1(n1568), .Y(n1101) );
  OAI222XL U2198 ( .A0(n1737), .A1(n1681), .B0(n2331), .B1(n1735), .C0(n1739), 
        .C1(n1490), .Y(n1100) );
  OAI222XL U2199 ( .A0(n1735), .A1(n1568), .B0(n1737), .B1(n1490), .C0(n1739), 
        .C1(n1681), .Y(n1099) );
  XNOR2X1 U2200 ( .A(n2541), .B(n2332), .Y(n1098) );
  XNOR2X1 U2201 ( .A(n1634), .B(n2333), .Y(n1096) );
  NOR2X1 U2202 ( .A(n2332), .B(n2334), .Y(n2333) );
  OAI22XL U2203 ( .A0(n2334), .A1(n2335), .B0(n2537), .B1(n2336), .Y(n1095) );
  OAI22XL U2204 ( .A0(n2335), .A1(n1792), .B0(n2538), .B1(n2339), .Y(n1094) );
  OAI22XL U2205 ( .A0(n2340), .A1(n2335), .B0(n2540), .B1(n2341), .Y(n1093) );
  OR3X1 U2206 ( .A(n2335), .B(n2541), .C(n2539), .Y(n2344) );
  NAND2X1 U2207 ( .A(n2345), .B(n1634), .Y(n2335) );
  OAI21XL U2208 ( .A0(n2346), .A1(n2338), .B0(HC3[0]), .Y(n2343) );
  OAI22XL U2209 ( .A0(n2334), .A1(n2347), .B0(n2534), .B1(n2348), .Y(n1091) );
  NAND2X1 U2210 ( .A(n2541), .B(n2539), .Y(n2334) );
  OAI22XL U2211 ( .A0(n1792), .A1(n2347), .B0(n2535), .B1(n2350), .Y(n1090) );
  NAND2X1 U2212 ( .A(n2539), .B(n1629), .Y(n1792) );
  OAI22XL U2213 ( .A0(n2340), .A1(n2347), .B0(n2536), .B1(n2351), .Y(n1089) );
  CLKINVX1 U2214 ( .A(n1793), .Y(n2340) );
  NOR2X1 U2215 ( .A(n1629), .B(n2539), .Y(n1793) );
  OAI31XL U2216 ( .A0(n2347), .A1(n2539), .A2(n2541), .B0(n2352), .Y(n1088) );
  OAI21XL U2217 ( .A0(n2346), .A1(n2349), .B0(HC3[4]), .Y(n2352) );
  OA21XL U2218 ( .A0(n2541), .A1(n2539), .B0(n2337), .Y(n2346) );
  NAND2X1 U2219 ( .A(n2542), .B(n2345), .Y(n2347) );
  AO22X1 U2220 ( .A0(n2353), .A1(n2354), .B0(n2355), .B1(n1711), .Y(n2345) );
  OAI22XL U2221 ( .A0(n1730), .A1(n1490), .B0(n1729), .B1(n1549), .Y(n2355) );
  OAI22XL U2222 ( .A0(n2609), .A1(n1728), .B0(n2583), .B1(n1828), .Y(n2353) );
  NAND2X1 U2223 ( .A(n799), .B(n2332), .Y(n1087) );
  OAI22XL U2224 ( .A0(n798), .A1(n1711), .B0(n799), .B1(n2356), .Y(n1086) );
  OAI22XL U2225 ( .A0(n797), .A1(n1711), .B0(n798), .B1(n2356), .Y(n1085) );
  OAI22XL U2226 ( .A0(n796), .A1(n1711), .B0(n797), .B1(n2356), .Y(n1084) );
  OAI22XL U2227 ( .A0(n795), .A1(n1711), .B0(n796), .B1(n2356), .Y(n1083) );
  OAI22XL U2228 ( .A0(n794), .A1(n1711), .B0(n795), .B1(n2356), .Y(n1082) );
  OAI22XL U2229 ( .A0(n793), .A1(n1711), .B0(n794), .B1(n2356), .Y(n1081) );
  OAI22XL U2230 ( .A0(n792), .A1(n1711), .B0(n793), .B1(n2356), .Y(n1080) );
  NAND2X1 U2231 ( .A(n2252), .B(n1711), .Y(n2356) );
  NOR2X1 U2232 ( .A(n2354), .B(n2342), .Y(n2332) );
  NOR2X1 U2233 ( .A(n2603), .B(n2609), .Y(n2326) );
  NOR2X1 U2234 ( .A(n2590), .B(n2596), .Y(n2329) );
  OAI21XL U2235 ( .A0(n2568), .A1(n2567), .B0(n2259), .Y(n2357) );
  NOR2X1 U2236 ( .A(n2577), .B(n2583), .Y(n2331) );
  OAI222XL U2237 ( .A0(n2154), .A1(n1664), .B0(n2359), .B1(n2184), .C0(n1714), 
        .C1(n1550), .Y(n1079) );
  OAI221XL U2238 ( .A0(n2146), .A1(n1514), .B0(n1713), .B1(n1664), .C0(n2360), 
        .Y(n1078) );
  AOI2BB2X1 U2239 ( .B0(n2149), .B1(n2616), .A0N(n1550), .A1N(n2150), .Y(n2360) );
  OAI221XL U2240 ( .A0(n1716), .A1(n1644), .B0(n1508), .B1(n1715), .C0(n2361), 
        .Y(n1077) );
  AOI2BB2X1 U2241 ( .B0(n2597), .B1(n2159), .A0N(n1717), .A1N(n1514), .Y(n2361) );
  OAI222XL U2242 ( .A0(n1562), .A1(n1718), .B0(n2162), .B1(n1514), .C0(n1719), 
        .C1(n1644), .Y(n1076) );
  OAI222XL U2243 ( .A0(n2188), .A1(n1501), .B0(n2362), .B1(n1720), .C0(n1721), 
        .C1(n1676), .Y(n1075) );
  OAI221XL U2244 ( .A0(n2189), .A1(n1676), .B0(n1723), .B1(n1514), .C0(n2363), 
        .Y(n1074) );
  OA22X1 U2245 ( .A0(n1722), .A1(n1569), .B0(n1724), .B1(n1501), .Y(n2363) );
  OAI222XL U2246 ( .A0(n1725), .A1(n1644), .B0(n2195), .B1(n1501), .C0(n1726), 
        .C1(n1569), .Y(n1073) );
  OAI222XL U2247 ( .A0(n1737), .A1(n1682), .B0(n2364), .B1(n1735), .C0(n1739), 
        .C1(n1491), .Y(n1072) );
  OAI222XL U2248 ( .A0(n1736), .A1(n1569), .B0(n1737), .B1(n1491), .C0(n1739), 
        .C1(n1682), .Y(n1071) );
  XNOR2X1 U2249 ( .A(n2550), .B(n2365), .Y(n1070) );
  XNOR2X1 U2250 ( .A(n1635), .B(n2366), .Y(n1068) );
  NOR2X1 U2251 ( .A(n2365), .B(n2367), .Y(n2366) );
  OAI22XL U2252 ( .A0(n2367), .A1(n2368), .B0(n2546), .B1(n2369), .Y(n1067) );
  OAI22XL U2253 ( .A0(n2368), .A1(n1788), .B0(n2547), .B1(n2372), .Y(n1066) );
  OAI22XL U2254 ( .A0(n2373), .A1(n2368), .B0(n2549), .B1(n2374), .Y(n1065) );
  OR3X1 U2255 ( .A(n2368), .B(n2550), .C(n2548), .Y(n2377) );
  NAND2X1 U2256 ( .A(n2378), .B(n1635), .Y(n2368) );
  OAI21XL U2257 ( .A0(n2379), .A1(n2371), .B0(HC2[0]), .Y(n2376) );
  OAI22XL U2258 ( .A0(n2367), .A1(n2380), .B0(n2543), .B1(n2381), .Y(n1063) );
  NAND2X1 U2259 ( .A(n2550), .B(n2548), .Y(n2367) );
  OAI22XL U2260 ( .A0(n1788), .A1(n2380), .B0(n2544), .B1(n2383), .Y(n1062) );
  NAND2X1 U2261 ( .A(n2548), .B(n1630), .Y(n1788) );
  OAI22XL U2262 ( .A0(n2373), .A1(n2380), .B0(n2545), .B1(n2384), .Y(n1061) );
  CLKINVX1 U2263 ( .A(n1789), .Y(n2373) );
  NOR2X1 U2264 ( .A(n1630), .B(n2548), .Y(n1789) );
  OAI31XL U2265 ( .A0(n2380), .A1(n2548), .A2(n2550), .B0(n2385), .Y(n1060) );
  OAI21XL U2266 ( .A0(n2379), .A1(n2382), .B0(HC2[4]), .Y(n2385) );
  OA21XL U2267 ( .A0(n2550), .A1(n2548), .B0(n2370), .Y(n2379) );
  NAND2X1 U2268 ( .A(n2551), .B(n2378), .Y(n2380) );
  AO22X1 U2269 ( .A0(n2386), .A1(n2387), .B0(n2388), .B1(n1712), .Y(n2378) );
  OAI22XL U2270 ( .A0(n1730), .A1(n1491), .B0(n1729), .B1(n1550), .Y(n2388) );
  OAI22XL U2271 ( .A0(n2610), .A1(n1728), .B0(n2584), .B1(n1828), .Y(n2386) );
  NAND2X1 U2272 ( .A(n778), .B(n2365), .Y(n1059) );
  OAI22XL U2273 ( .A0(n777), .A1(n1712), .B0(n778), .B1(n2389), .Y(n1058) );
  OAI22XL U2274 ( .A0(n776), .A1(n1712), .B0(n777), .B1(n2389), .Y(n1057) );
  OAI22XL U2275 ( .A0(n775), .A1(n1712), .B0(n776), .B1(n2389), .Y(n1056) );
  OAI22XL U2276 ( .A0(n774), .A1(n1712), .B0(n775), .B1(n2389), .Y(n1055) );
  OAI22XL U2277 ( .A0(n773), .A1(n1712), .B0(n774), .B1(n2389), .Y(n1054) );
  OAI22XL U2278 ( .A0(n772), .A1(n1712), .B0(n773), .B1(n2389), .Y(n1053) );
  OAI22XL U2279 ( .A0(n771), .A1(n1712), .B0(n772), .B1(n2389), .Y(n1052) );
  NAND2X1 U2280 ( .A(n2252), .B(n1712), .Y(n2389) );
  NOR2X1 U2281 ( .A(n2387), .B(n2375), .Y(n2365) );
  OAI211X1 U2282 ( .A0(n2364), .A1(n2254), .B0(n2390), .C0(n2391), .Y(n2387)
         );
  NOR2X1 U2283 ( .A(n2604), .B(n2610), .Y(n2359) );
  NOR2X1 U2284 ( .A(n2591), .B(n2597), .Y(n2362) );
  OAI21XL U2285 ( .A0(n2570), .A1(n2569), .B0(n2259), .Y(n2390) );
  NOR2X1 U2286 ( .A(n2578), .B(n2584), .Y(n2364) );
  OAI222XL U2287 ( .A0(n2154), .A1(n1665), .B0(n2392), .B1(n2184), .C0(n1714), 
        .C1(n1551), .Y(n1051) );
  NAND2X1 U2288 ( .A(n1614), .B(n1714), .Y(n2184) );
  OAI221XL U2289 ( .A0(n2146), .A1(n1515), .B0(n1713), .B1(n1665), .C0(n2393), 
        .Y(n1050) );
  AOI2BB2X1 U2290 ( .B0(n2149), .B1(n2617), .A0N(n1551), .A1N(n2150), .Y(n2393) );
  OA22X1 U2291 ( .A0(\C2[2][7] ), .A1(n942), .B0(n2397), .B1(n2398), .Y(n2396)
         );
  NOR2BX1 U2292 ( .AN(n942), .B(n943), .Y(n2398) );
  AOI32X1 U2293 ( .A0(n2399), .A1(n2400), .A2(n2401), .B0(n2402), .B1(n2403), 
        .Y(n2397) );
  OAI21XL U2294 ( .A0(n2404), .A1(n937), .B0(\C2[2][6] ), .Y(n2403) );
  NAND2X1 U2295 ( .A(n2404), .B(n937), .Y(n2402) );
  AOI32X1 U2296 ( .A0(n930), .A1(\C2[3][4] ), .A2(n2400), .B0(\C2[3][5] ), 
        .B1(n934), .Y(n2404) );
  AOI2BB2X1 U2297 ( .B0(n937), .B1(\C2[2][6] ), .A0N(n930), .A1N(\C2[3][4] ), 
        .Y(n2401) );
  NAND2X1 U2298 ( .A(n933), .B(\C2[2][5] ), .Y(n2400) );
  OAI211X1 U2299 ( .A0(n925), .A1(n2405), .B0(n2406), .C0(n2407), .Y(n2399) );
  AO21X1 U2300 ( .A0(n2405), .A1(n925), .B0(\C2[2][3] ), .Y(n2407) );
  OAI222XL U2301 ( .A0(n926), .A1(\C2[3][3] ), .B0(n922), .B1(\C2[3][2] ), 
        .C0(n2408), .C1(n2409), .Y(n2406) );
  NOR2X1 U2302 ( .A(n917), .B(\C2[2][1] ), .Y(n2409) );
  AOI211X1 U2303 ( .A0(n917), .A1(\C2[2][1] ), .B0(\C2[2][0] ), .C0(n945), .Y(
        n2408) );
  NAND2X1 U2304 ( .A(n922), .B(\C2[3][2] ), .Y(n2405) );
  CLKINVX1 U2305 ( .A(n1845), .Y(n1838) );
  OAI221XL U2306 ( .A0(n1716), .A1(n1645), .B0(n1509), .B1(n1715), .C0(n2410), 
        .Y(n1049) );
  AOI2BB2X1 U2307 ( .B0(n2598), .B1(n2159), .A0N(n1717), .A1N(n1515), .Y(n2410) );
  CLKINVX1 U2308 ( .A(n2394), .Y(n2395) );
  OAI22XL U2309 ( .A0(n943), .A1(n1607), .B0(n2412), .B1(n2413), .Y(n2411) );
  NOR2X1 U2310 ( .A(n941), .B(\C2[2][7] ), .Y(n2413) );
  AOI32X1 U2311 ( .A0(n2414), .A1(n2415), .A2(n2416), .B0(n2417), .B1(n2418), 
        .Y(n2412) );
  OAI21XL U2312 ( .A0(n2419), .A1(n1617), .B0(n938), .Y(n2418) );
  NAND2X1 U2313 ( .A(n2419), .B(n1617), .Y(n2417) );
  AOI32X1 U2314 ( .A0(n928), .A1(\C2[2][4] ), .A2(n2415), .B0(\C2[2][5] ), 
        .B1(n932), .Y(n2419) );
  AOI2BB2X1 U2315 ( .B0(n1532), .B1(n930), .A0N(\C2[2][6] ), .A1N(n936), .Y(
        n2416) );
  NAND2X1 U2316 ( .A(n934), .B(n1585), .Y(n2415) );
  OAI211X1 U2317 ( .A0(n926), .A1(n2420), .B0(n2421), .C0(n2422), .Y(n2414) );
  AO21X1 U2318 ( .A0(n2420), .A1(n926), .B0(n1601), .Y(n2422) );
  OAI222XL U2319 ( .A0(n924), .A1(\C2[2][3] ), .B0(n920), .B1(\C2[2][2] ), 
        .C0(n2423), .C1(n2424), .Y(n2421) );
  AND2X1 U2320 ( .A(n916), .B(\C2[2][1] ), .Y(n2424) );
  CLKINVX1 U2321 ( .A(n2425), .Y(n2423) );
  OAI211X1 U2322 ( .A0(\C2[2][1] ), .A1(n916), .B0(n944), .C0(\C2[2][0] ), .Y(
        n2425) );
  NAND2X1 U2323 ( .A(n920), .B(\C2[2][2] ), .Y(n2420) );
  OAI222XL U2324 ( .A0(n1563), .A1(n1718), .B0(n2162), .B1(n1515), .C0(n1719), 
        .C1(n1645), .Y(n1048) );
  AOI2BB2X1 U2325 ( .B0(n940), .B1(n1607), .A0N(n2427), .A1N(n2428), .Y(n2426)
         );
  NOR2X1 U2326 ( .A(n940), .B(n1607), .Y(n2428) );
  AOI32X1 U2327 ( .A0(n2429), .A1(n2430), .A2(n2431), .B0(n2432), .B1(n2433), 
        .Y(n2427) );
  OAI21XL U2328 ( .A0(n2434), .A1(n1595), .B0(n936), .Y(n2433) );
  NAND2X1 U2329 ( .A(n2434), .B(n1595), .Y(n2432) );
  AOI32X1 U2330 ( .A0(n927), .A1(n1532), .A2(n2430), .B0(n1585), .B1(n931), 
        .Y(n2434) );
  AOI2BB2X1 U2331 ( .B0(n936), .B1(n1595), .A0N(n1532), .A1N(n927), .Y(n2431)
         );
  OR2X1 U2332 ( .A(n931), .B(n1585), .Y(n2430) );
  OAI211X1 U2333 ( .A0(n924), .A1(n2435), .B0(n2436), .C0(n2437), .Y(n2429) );
  OAI2BB1X1 U2334 ( .A0N(n2435), .A1N(n924), .B0(n923), .Y(n2437) );
  OAI222XL U2335 ( .A0(n923), .A1(n1601), .B0(n919), .B1(n1534), .C0(n2438), 
        .C1(n2439), .Y(n2436) );
  NOR2X1 U2336 ( .A(n916), .B(n1537), .Y(n2439) );
  AOI211X1 U2337 ( .A0(n916), .A1(n1537), .B0(n1603), .C0(n944), .Y(n2438) );
  NAND2X1 U2338 ( .A(n919), .B(n1534), .Y(n2435) );
  CLKINVX1 U2339 ( .A(n1842), .Y(n2102) );
  NOR3X1 U2340 ( .A(sort_stage[0]), .B(sort_stage[2]), .C(n1581), .Y(n1842) );
  OAI222XL U2341 ( .A0(n2188), .A1(n1502), .B0(n2440), .B1(n1720), .C0(n1721), 
        .C1(n1677), .Y(n1047) );
  OAI221XL U2342 ( .A0(n2189), .A1(n1677), .B0(n1723), .B1(n1515), .C0(n2442), 
        .Y(n1046) );
  OA22X1 U2343 ( .A0(n1722), .A1(n1570), .B0(n1724), .B1(n1502), .Y(n2442) );
  NAND3X1 U2344 ( .A(n1844), .B(n2443), .C(n1845), .Y(n2441) );
  OAI22XL U2345 ( .A0(n914), .A1(\C3[1][7] ), .B0(n2444), .B1(n2445), .Y(n2443) );
  NOR2BX1 U2346 ( .AN(n914), .B(n913), .Y(n2445) );
  AOI32X1 U2347 ( .A0(n2446), .A1(n2447), .A2(n2448), .B0(n2449), .B1(n2450), 
        .Y(n2444) );
  OAI21XL U2348 ( .A0(n2451), .A1(\C3[1][6] ), .B0(n893), .Y(n2450) );
  NAND2X1 U2349 ( .A(n2451), .B(\C3[1][6] ), .Y(n2449) );
  CLKINVX1 U2350 ( .A(n2452), .Y(n2451) );
  OAI32X1 U2351 ( .A0(\C3[1][4] ), .A1(n899), .A2(n2453), .B0(n896), .B1(
        \C3[1][5] ), .Y(n2452) );
  CLKINVX1 U2352 ( .A(n2447), .Y(n2453) );
  AOI22X1 U2353 ( .A0(\C3[1][6] ), .A1(n893), .B0(n899), .B1(\C3[1][4] ), .Y(
        n2448) );
  NAND2X1 U2354 ( .A(n896), .B(\C3[1][5] ), .Y(n2447) );
  OAI211X1 U2355 ( .A0(n902), .A1(n2454), .B0(n2455), .C0(n2456), .Y(n2446) );
  AO21X1 U2356 ( .A0(n2454), .A1(n902), .B0(\C3[1][3] ), .Y(n2456) );
  OAI222XL U2357 ( .A0(n904), .A1(\C3[2][2] ), .B0(n901), .B1(\C3[2][3] ), 
        .C0(n2457), .C1(n2458), .Y(n2455) );
  NOR2X1 U2358 ( .A(n908), .B(\C3[1][1] ), .Y(n2458) );
  AOI211X1 U2359 ( .A0(n908), .A1(\C3[1][1] ), .B0(\C3[1][0] ), .C0(n910), .Y(
        n2457) );
  NAND2X1 U2360 ( .A(n904), .B(\C3[2][2] ), .Y(n2454) );
  OAI222XL U2361 ( .A0(n1725), .A1(n1645), .B0(n2195), .B1(n1502), .C0(n1726), 
        .C1(n1570), .Y(n1045) );
  AOI2BB2X1 U2362 ( .B0(n912), .B1(\C3[1][7] ), .A0N(n2460), .A1N(n2461), .Y(
        n2459) );
  NOR2X1 U2363 ( .A(n912), .B(\C3[1][7] ), .Y(n2461) );
  AOI32X1 U2364 ( .A0(n2462), .A1(n2463), .A2(n2464), .B0(n2465), .B1(n2466), 
        .Y(n2460) );
  OAI21XL U2365 ( .A0(n2467), .A1(n1599), .B0(n892), .Y(n2466) );
  NAND2X1 U2366 ( .A(n2467), .B(n1599), .Y(n2465) );
  AOI32X1 U2367 ( .A0(n897), .A1(\C3[1][4] ), .A2(n2463), .B0(\C3[1][5] ), 
        .B1(n894), .Y(n2467) );
  OA22X1 U2368 ( .A0(\C3[1][6] ), .A1(n891), .B0(\C3[1][4] ), .B1(n897), .Y(
        n2464) );
  OR2X1 U2369 ( .A(n894), .B(\C3[1][5] ), .Y(n2463) );
  OAI211X1 U2370 ( .A0(n901), .A1(n2468), .B0(n2469), .C0(n2470), .Y(n2462) );
  OAI2BB1X1 U2371 ( .A0N(n2468), .A1N(n901), .B0(n900), .Y(n2470) );
  OAI222XL U2372 ( .A0(n903), .A1(\C3[1][2] ), .B0(n900), .B1(\C3[1][3] ), 
        .C0(n2471), .C1(n2472), .Y(n2469) );
  AND2X1 U2373 ( .A(n906), .B(\C3[1][1] ), .Y(n2472) );
  CLKINVX1 U2374 ( .A(n2473), .Y(n2471) );
  OAI211X1 U2375 ( .A0(\C3[1][1] ), .A1(n906), .B0(n909), .C0(\C3[1][0] ), .Y(
        n2473) );
  NAND2X1 U2376 ( .A(n903), .B(\C3[1][2] ), .Y(n2468) );
  OAI222XL U2377 ( .A0(n1737), .A1(n1683), .B0(n2474), .B1(n1735), .C0(n1739), 
        .C1(n1492), .Y(n1044) );
  OAI222XL U2378 ( .A0(n1736), .A1(n1570), .B0(n1737), .B1(n1492), .C0(n1739), 
        .C1(n1683), .Y(n1043) );
  NAND3X1 U2379 ( .A(n1845), .B(n1846), .C(N2784), .Y(n2475) );
  NOR3X1 U2380 ( .A(sort_stage[1]), .B(sort_stage[2]), .C(sort_stage[0]), .Y(
        n1845) );
  XNOR2X1 U2381 ( .A(n2559), .B(n2476), .Y(n1042) );
  XNOR2X1 U2382 ( .A(n1636), .B(n2477), .Y(n1040) );
  NOR2X1 U2383 ( .A(n2476), .B(n2478), .Y(n2477) );
  NAND2X1 U2384 ( .A(n758), .B(n2476), .Y(n1039) );
  OAI22XL U2385 ( .A0(n757), .A1(n1727), .B0(n758), .B1(n2479), .Y(n1038) );
  OAI22XL U2386 ( .A0(n756), .A1(n1727), .B0(n757), .B1(n2479), .Y(n1037) );
  OAI22XL U2387 ( .A0(n755), .A1(n1727), .B0(n756), .B1(n2479), .Y(n1036) );
  OAI22XL U2388 ( .A0(n754), .A1(n1727), .B0(n755), .B1(n2479), .Y(n1035) );
  OAI22XL U2389 ( .A0(n753), .A1(n1727), .B0(n754), .B1(n2479), .Y(n1034) );
  OAI22XL U2390 ( .A0(n752), .A1(n1727), .B0(n753), .B1(n2479), .Y(n1033) );
  OAI22XL U2391 ( .A0(n751), .A1(n1727), .B0(n752), .B1(n2479), .Y(n1032) );
  NAND2X1 U2392 ( .A(n1727), .B(n2252), .Y(n2479) );
  NAND3X1 U2393 ( .A(n1730), .B(n1729), .C(n1820), .Y(n2252) );
  NOR2X1 U2394 ( .A(n1824), .B(n1846), .Y(n1820) );
  OAI22XL U2395 ( .A0(n2478), .A1(n2480), .B0(n2552), .B1(n2481), .Y(n1031) );
  OAI22XL U2396 ( .A0(n2480), .A1(n1784), .B0(n2553), .B1(n2484), .Y(n1030) );
  OAI22XL U2397 ( .A0(n2485), .A1(n2480), .B0(n2554), .B1(n2486), .Y(n1029) );
  OAI31XL U2398 ( .A0(n2480), .A1(n2557), .A2(n2559), .B0(n2488), .Y(n1028) );
  OAI21XL U2399 ( .A0(n2489), .A1(n2483), .B0(HC1[4]), .Y(n2488) );
  NAND2X1 U2400 ( .A(n2560), .B(n2490), .Y(n2480) );
  OAI22XL U2401 ( .A0(n2478), .A1(n2491), .B0(n2555), .B1(n2492), .Y(n1027) );
  NAND2X1 U2402 ( .A(n2559), .B(n2557), .Y(n2478) );
  OAI22XL U2403 ( .A0(n1784), .A1(n2491), .B0(n2556), .B1(n2494), .Y(n1026) );
  NAND2X1 U2404 ( .A(n2557), .B(n1631), .Y(n1784) );
  OAI22XL U2405 ( .A0(n2485), .A1(n2491), .B0(n2558), .B1(n2495), .Y(n1025) );
  CLKINVX1 U2406 ( .A(n1785), .Y(n2485) );
  NOR2X1 U2407 ( .A(n1631), .B(n2557), .Y(n1785) );
  OR3X1 U2408 ( .A(n2491), .B(n2559), .C(n2557), .Y(n2497) );
  NAND2X1 U2409 ( .A(n2490), .B(n1636), .Y(n2491) );
  AO22X1 U2410 ( .A0(n2498), .A1(n2499), .B0(n2500), .B1(n1727), .Y(n2490) );
  OAI22XL U2411 ( .A0(n1730), .A1(n1492), .B0(n1729), .B1(n1551), .Y(n2500) );
  OAI22XL U2412 ( .A0(n2611), .A1(n1728), .B0(n2585), .B1(n1828), .Y(n2498) );
  OAI21XL U2413 ( .A0(n2489), .A1(n2493), .B0(HC1[0]), .Y(n2496) );
  NOR2X1 U2414 ( .A(n2499), .B(n2487), .Y(n2476) );
  OAI211X1 U2415 ( .A0(n2474), .A1(n2254), .B0(n2501), .C0(n2502), .Y(n2499)
         );
  NOR2X1 U2416 ( .A(n2605), .B(n2611), .Y(n2392) );
  CLKINVX1 U2417 ( .A(n1728), .Y(n1824) );
  NOR3X1 U2418 ( .A(state[0]), .B(state[2]), .C(gray_valid), .Y(n1994) );
  NOR2X1 U2419 ( .A(n2592), .B(n2598), .Y(n2440) );
  CLKINVX1 U2420 ( .A(n1729), .Y(n1844) );
  OAI21XL U2421 ( .A0(n2572), .A1(n2571), .B0(n2259), .Y(n2501) );
  CLKINVX1 U2422 ( .A(n1730), .Y(n2259) );
  NAND2X1 U2423 ( .A(n1846), .B(n1613), .Y(n2254) );
  NOR3X1 U2424 ( .A(gray_valid), .B(state[1]), .C(n1586), .Y(n2504) );
  NOR2X1 U2425 ( .A(n2579), .B(n2585), .Y(n2474) );
  OA21XL U2426 ( .A0(n2559), .A1(n2557), .B0(n2482), .Y(n2489) );
  NAND2X1 U2427 ( .A(n2503), .B(n1583), .Y(n1822) );
  NOR3X1 U2428 ( .A(gray_valid), .B(state[2]), .C(n1580), .Y(n2503) );
endmodule

